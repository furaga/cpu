library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
entity fadd is
	port (
		I1, I2 : in  std_logic_vector (0 to 31);
		O  : out std_logic_vector (0 to 31));
end fadd;

architecture fadd_archi of fadd is

	signal s1, s2 : std_logic;
	signal e1, e2 : std_logic_vector(0 to 7);
	signal c1, c2 : std_logic_vector(0 to 23);
	signal E1I, E2I, C1I, C2I : integer;

begin  -- fadd_archi

	s1 <= I1(0);
	s2 <= I2(0);
	e1(0 to 7) <= I1(1 to 8);
	e2(0 to 7) <= I2(1 to 8);
	c1(0 to 23) <= '1'&I1(9 to 31);
	c2(0 to 23) <= '1'&I2(9 to 31);

	E1I <= conv_integer(e1(0 to 7));
	E2I <= conv_integer(e2(0 to 7));
	C1I <= conv_integer(c1(0 to 23));
	C2I <= conv_integer(c2(0 to 23));
  
  	add :process(I1,I2)
		variable S3 : std_logic := '0';
		variable E3V : std_logic_vector(0 to 7);
		variable E3VI : integer;
		variable C1V, C2V : std_logic_vector(0 to 23);
		variable C3V : std_logic_vector(0 to 24);
		variable C3VA : std_logic_vector(0 to 24) := conv_std_logic_vector(0, 25);
		variable COUNT : integer := 25;
		
	  begin
		if true then
			if E1I=0 then 
				O <= I2;
			elsif E2I=0 then 
				O <= I1;
			else 
				O <= x"12345678";
			end if;
		else


      if (S1 = '1' and S2 = '1') or ((S1 = '1') and ((E1I > E2I) or ((E1I = E2I) and (C1I > C2I)))) or ((S2 = '1') and ((E1I < E2I) or ((E1I = E2I) and (C1I < C2I)))) then
        S3 := '1';
      else s3 := '0';
      end if;
    
      if E1I < E2I then
        E3V := E2;
        if (E2I - E1I) < 24 then
          C1V((E2I - E1I) to 23) := C1(0 to (23 - (E2I - E1I)));
          C1V(0 to (E2I - E1I -1)) := C1(0 to (E2I - E1I - 1)) - C1(0 to (E2I - E1I - 1));
        else
          C1V := conv_std_logic_vector(0, 24);
        end if;
        C2V := C2;
      
      else
        E3V := E1;
        if (E1I - E2I) < 24 then
          C2V((E1I - E2I) to 23)  := C2(0 to (23 - (E1I - E2I)));
          C2V(0 to (E1I - E2I -1)) := C2(0 to (E1I - E2I - 1)) - C2(0 to (E1I - E2I - 1));
        else
          C2V := conv_std_logic_vector(0, 24);
        end if;
        C1V := C1;          
      end if;
    
      E3VI := conv_integer(E3V);
    
      if S1 = S2 then
        C3V(0 to 24) := ('0' & C1V(0 to 23)) + ('0' & C2V(0 to 23));
      else
        if C1V > C2V then
          C3V(0 to 24) := ('0' & C1V(0 to 23)) - ('0' & C2V(0 to 23));
        else
          C3V(0 to 24) := ('0' & C2V(0 to 23)) - ('0' & C1V(0 to 23));
        end if;
      end if;
    
      for I in C3V'range loop
        if C3V(I) = '1' then
          if COUNT = 25  then
            COUNT := I;
          end if;
        end if;
      end loop;
    
      C3VA := conv_std_logic_vector(0, 25);
      E3VI := E3VI - COUNT + 1;
      E3V := conv_std_logic_vector(E3VI, 8);
      if COUNT = 0 then
        C3VA(1 to 24) := C3V(0 to 23);
      elsif COUNT = 25 then
        E3V := conv_std_logic_vector(0, 8);
      else
        C3VA(1 to (25 - COUNT)) := C3V(COUNT to 24);
      end if;
      COUNT := 25;
      O <= S3 & E3V & C3VA(2 to 24);


	end if;

  end process;

end fadd_archi;
