library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is
	port (
		clka : in std_logic;
		addra : in std_logic_vector(13 downto 0);
		douta : out std_logic_vector(31 downto 0));



end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 32767) of word_t;
	signal addr_in	: integer range 0 to 32767;

	constant mem : mem_t := (
x"000000F4",
x"00000000",
x"3F800000",
x"BF800000",
x"00800000",
x"4B000000",
x"4B000000",
x"43160000",
x"C3160000",
x"C0000000",
x"3B800000",
x"41A00000",
x"3D4CCCC4",
x"3E800000",
x"41200000",
x"3E999999",
x"3E199999",
x"40490FDA",
x"41F00000",
x"BFC90FDA",
x"40800000",
x"41800000",
x"41300000",
x"41C80000",
x"41500000",
x"42100000",
x"42440000",
x"41880000",
x"42800000",
x"41980000",
x"42A20000",
x"41A80000",
x"42C80000",
x"41B80000",
x"42F20000",
x"41700000",
x"38D1B70F",
x"4CBEBC20",
x"BDCCCCC4",
x"3C23D70A",
x"BE4CCCC4",
x"BF800000",
x"3DCCCCC4",
x"3F66665E",
x"3E4CCCC4",
x"C3480000",
x"43480000",
x"40400000",
x"40A00000",
x"41100000",
x"40E00000",
x"3F800000",
x"3C8EFA2D",
x"43000000",
x"4E6E6B28",
x"437F0000",
x"00000000",
x"3FC90FDA",
x"3F000000",
x"40C90FDA",
x"40000000",
x"40490FDA",
x"080000D3",
x"A0630002",
x"00622820",
x"20430000",
x"68A20005",
x"28A20004",
x"AC440000",
x"20420004",
x"08000042",
x"E0000000",
x"A0630002",
x"00622020",
x"20430000",
x"68820005",
x"28820004",
x"E4400000",
x"20420004",
x"0800004B",
x"E0000000",
x"44000806",
x"20030000",
x"C4640000",
x"E8800015",
x"C8800014",
x"44000007",
x"20030010",
x"C4620000",
x"E8020004",
x"C8020003",
x"44000007",
x"E0000000",
x"44020000",
x"44020001",
x"44200807",
x"E820001B",
x"C820001A",
x"44020000",
x"20030004",
x"C4630000",
x"44030000",
x"44020001",
x"44000007",
x"E0000000",
x"20030010",
x"C4620000",
x"E8020003",
x"C8020002",
x"E0000000",
x"44000806",
x"44020000",
x"E4200000",
x"8C240000",
x"44020001",
x"E4200000",
x"8C240000",
x"E8010005",
x"C8010004",
x"20030004",
x"C4630000",
x"44030001",
x"E0000000",
x"44000007",
x"E0000000",
x"44000007",
x"C0000051",
x"44000007",
x"E0000000",
x"68030006",
x"28030005",
x"00031822",
x"C0000087",
x"44000007",
x"E0000000",
x"20050010",
x"C4A10000",
x"20050014",
x"8CA40000",
x"2005000C",
x"8CA50000",
x"68A30007",
x"28A30006",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"E0000000",
x"20040000",
x"C4820000",
x"00651822",
x"44411000",
x"68A3FFFE",
x"28A3FFFD",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"44020000",
x"E0000000",
x"20030000",
x"C4610000",
x"E8200006",
x"C8200005",
x"44000007",
x"C00000A8",
x"00031822",
x"E0000000",
x"C0000051",
x"20040010",
x"C4820000",
x"20040014",
x"8C840000",
x"E8400007",
x"C8400006",
x"44020000",
x"E4200000",
x"8C230000",
x"00641822",
x"E0000000",
x"2005000C",
x"8CA50000",
x"20030000",
x"44020001",
x"00651820",
x"E840FFFE",
x"C840FFFD",
x"44020000",
x"E4200000",
x"8C250000",
x"00A42822",
x"00A31820",
x"E0000000",
x"080000A0",
x"20030000",
x"04002000",
x"00641820",
x"A0630008",
x"04002000",
x"00641820",
x"A0630008",
x"04002000",
x"00641820",
x"A0630008",
x"04002000",
x"00641820",
x"E0000000",
x"C00000C2",
x"AC230000",
x"C4200000",
x"E0000000",
x"203F0000",
x"40210940",
x"201C0001",
x"201DFFFF",
x"201B00DC",
x"C7700000",
x"201B00C8",
x"C7710000",
x"201B0018",
x"C7720000",
x"201B001C",
x"C7730000",
x"201B00A0",
x"C7740000",
x"201B00E4",
x"C7750000",
x"201B00E0",
x"C7760000",
x"201B00B8",
x"C7770000",
x"201B00BC",
x"C7780000",
x"201B00C0",
x"C7790000",
x"201B00C4",
x"C77A0000",
x"201B00D8",
x"C77B0000",
x"201B0088",
x"C77C0000",
x"201B00E8",
x"C77D0000",
x"201B0040",
x"C77E0000",
x"201B0048",
x"C77F0000",
x"200300F0",
x"C4640000",
x"200300EC",
x"C46A0000",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20004",
x"40210004",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20008",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E2000C",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20010",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040001",
x"AFE2093C",
x"43E20014",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20018",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E2001C",
x"C000003F",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E20020",
x"46000006",
x"C0000048",
x"20640000",
x"8FE2093C",
x"2006003C",
x"200A0000",
x"20090000",
x"20080000",
x"20070000",
x"20050000",
x"20430000",
x"2042002C",
x"AC64FFD8",
x"AC64FFDC",
x"AC64FFE0",
x"AC64FFE4",
x"AC65FFE8",
x"AC64FFEC",
x"AC64FFF0",
x"AC67FFF4",
x"AC68FFF8",
x"AC69FFFC",
x"AC6A0000",
x"AFE2093C",
x"43E20110",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2011C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20128",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20134",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030001",
x"AFE2093C",
x"43E20138",
x"47600006",
x"C0000048",
x"8FE2093C",
x"20060032",
x"20030001",
x"2004FFFF",
x"C000003F",
x"20640000",
x"AFE2093C",
x"43E20200",
x"20C30000",
x"C000003F",
x"8FE2093C",
x"20060001",
x"20030001",
x"8FE40200",
x"C000003F",
x"20640000",
x"AFE2093C",
x"43E20204",
x"20C30000",
x"C000003F",
x"8FE2093C",
x"20030001",
x"AFE2093C",
x"43E20208",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E2020C",
x"C000003F",
x"8FE2093C",
x"20030001",
x"200400D4",
x"C4800000",
x"AFE2093C",
x"43E20210",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2021C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20220",
x"C000003F",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2022C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20238",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20244",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20250",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030002",
x"20040000",
x"AFE2093C",
x"43E20258",
x"C000003F",
x"8FE2093C",
x"20030002",
x"20040000",
x"AFE2093C",
x"43E20260",
x"C000003F",
x"8FE2093C",
x"20030001",
x"AFE2093C",
x"43E20264",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20270",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2027C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20288",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20294",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E202A0",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E202AC",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E202B0",
x"46000006",
x"C0000048",
x"20670000",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E202B4",
x"43E402B0",
x"C000003F",
x"20640000",
x"8FE2093C",
x"20060000",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"AFE2093C",
x"43E202B8",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E202CC",
x"43E402B8",
x"C000003F",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E202D0",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E202DC",
x"46000006",
x"C0000048",
x"20660000",
x"8FE2093C",
x"2003003C",
x"AFE2093C",
x"43E203CC",
x"43E402D0",
x"C000003F",
x"20640000",
x"8FE2093C",
x"AFE2093C",
x"43E203D4",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC660000",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E203D8",
x"46000006",
x"C0000048",
x"20660000",
x"8FE2093C",
x"20030000",
x"AFE2093C",
x"43E203DC",
x"43E403D8",
x"C000003F",
x"8FE2093C",
x"AFE2093C",
x"43E203E4",
x"20440000",
x"20420008",
x"AC83FFFC",
x"AC860000",
x"8FE2093C",
x"200600B4",
x"20050000",
x"20430000",
x"2042000C",
x"E470FFF8",
x"AC64FFFC",
x"AC650000",
x"AFE2093C",
x"43E206B4",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE2093C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E206B8",
x"C000003F",
x"8FE2093C",
x"20030080",
x"20040080",
x"AFE30258",
x"AFE40254",
x"20040040",
x"AFE40260",
x"20040040",
x"AFE4025C",
x"200400D0",
x"C4830000",
x"C0000081",
x"44600003",
x"E7E00264",
x"8FEC0258",
x"20030003",
x"AFE2093C",
x"43E206C4",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E206D0",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E206E4",
x"43E406D0",
x"C000003F",
x"206A0000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306E0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306DC",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306D8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306D4",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E206F8",
x"C000003F",
x"20690000",
x"8FE2093C",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E2070C",
x"C000003F",
x"20680000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20718",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E2072C",
x"43E40718",
x"C000003F",
x"20670000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30728",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30724",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30720",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3071C",
x"20030003",
x"AFE2093C",
x"43E20738",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E2074C",
x"43E40738",
x"C000003F",
x"20660000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30748",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30744",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30740",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3073C",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20750",
x"C000003F",
x"206D0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2075C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E20770",
x"43E4075C",
x"C000003F",
x"20650000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3076C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30768",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30764",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30760",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA0774",
x"8FE30258",
x"40690002",
x"C0002F38",
x"20710000",
x"AFF10778",
x"8FEC0258",
x"20030003",
x"AFE2093C",
x"43E20784",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20790",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E207A4",
x"43E40790",
x"C000003F",
x"206A0000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307A0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3079C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30798",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30794",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E207B8",
x"C000003F",
x"20690000",
x"8FE2093C",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E207CC",
x"C000003F",
x"20680000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E207D8",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E207EC",
x"43E407D8",
x"C000003F",
x"20670000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307DC",
x"20030003",
x"AFE2093C",
x"43E207F8",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E2080C",
x"43E407F8",
x"C000003F",
x"20660000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30808",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30804",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30800",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307FC",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E20810",
x"C000003F",
x"206D0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E2081C",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E20830",
x"43E4081C",
x"C000003F",
x"20650000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3082C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30828",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30824",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30820",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA0834",
x"8FE30258",
x"40690002",
x"C0002F38",
x"20700000",
x"AFF00838",
x"8FEC0258",
x"20030003",
x"AFE2093C",
x"43E20844",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20850",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E20864",
x"43E40850",
x"C000003F",
x"206A0000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30860",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3085C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30858",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30854",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E20878",
x"C000003F",
x"20690000",
x"8FE2093C",
x"20030005",
x"20040000",
x"AFE2093C",
x"43E2088C",
x"C000003F",
x"20680000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E20898",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E208AC",
x"43E40898",
x"C000003F",
x"20670000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3089C",
x"20030003",
x"AFE2093C",
x"43E208B8",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E208CC",
x"43E408B8",
x"C000003F",
x"20660000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308BC",
x"20030001",
x"20040000",
x"AFE2093C",
x"43E208D0",
x"C000003F",
x"206D0000",
x"8FE2093C",
x"20030003",
x"AFE2093C",
x"43E208DC",
x"46000006",
x"C0000048",
x"8FE2093C",
x"20030005",
x"AFE2093C",
x"43E208F0",
x"43E408DC",
x"C000003F",
x"20650000",
x"8FE2093C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308EC",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E0",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA08F4",
x"8FE30258",
x"40690002",
x"C0002F38",
x"20210004",
x"206F0000",
x"AFEF08F8",
x"AC310000",
x"AC2F0004",
x"AC300008",
x"E42A000C",
x"E4240010",
x"40210018",
x"C00000CF",
x"E7E0011C",
x"C00000CF",
x"E7E00118",
x"C00000CF",
x"E7E00114",
x"C00000CF",
x"20210018",
x"200300CC",
x"C4670000",
x"44071802",
x"46C31001",
x"E8500003",
x"44400806",
x"08000453",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000479",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800046A",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000465",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"0800046A",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"08000479",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000474",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"08000479",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"0800049C",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800048D",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000488",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"0800048D",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"0800049C",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000497",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"0800049C",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"C4240010",
x"E8800006",
x"EA020003",
x"20030000",
x"080004A2",
x"20030001",
x"080004A7",
x"EA020003",
x"20030001",
x"080004A7",
x"20030000",
x"E8800003",
x"44000806",
x"080004AB",
x"47A00801",
x"EAC10003",
x"44200006",
x"080004AF",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"C42A000C",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44003007",
x"080004C3",
x"44003006",
x"E8700003",
x"44600806",
x"080004C7",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080004ED",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080004DE",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080004D9",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"080004DE",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"080004ED",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080004E8",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"080004ED",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"08000510",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000501",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080004FC",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"08000501",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"08000510",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800050B",
x"443D0800",
x"40210018",
x"C0000A77",
x"20210018",
x"08000510",
x"443D0801",
x"40210018",
x"C0000A77",
x"20210018",
x"E8800006",
x"EA030003",
x"20030000",
x"08000515",
x"20030001",
x"0800051A",
x"EA030003",
x"20030001",
x"0800051A",
x"20030000",
x"E8800003",
x"44000806",
x"0800051E",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000522",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44002807",
x"08000535",
x"44002806",
x"E4250014",
x"E4260018",
x"E427001C",
x"40210024",
x"C00000CF",
x"20210024",
x"C427001C",
x"44071802",
x"46C31001",
x"E8500003",
x"44400806",
x"08000542",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000568",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000559",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000554",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"08000559",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"08000568",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000563",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"08000568",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"0800058B",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800057C",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000577",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"0800057C",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"0800058B",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000586",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"0800058B",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"C4240010",
x"E8800006",
x"EA020003",
x"20030000",
x"08000591",
x"20030001",
x"08000596",
x"EA020003",
x"20030001",
x"08000596",
x"20030000",
x"E8800003",
x"44000806",
x"0800059A",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800059E",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"C42A000C",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44001007",
x"080005B2",
x"44001006",
x"E8700003",
x"44600806",
x"080005B6",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080005DC",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080005CD",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005C8",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"080005CD",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"080005DC",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005D7",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"080005DC",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"080005FF",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080005F0",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005EB",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"080005F0",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"080005FF",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005FA",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"080005FF",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"E8800006",
x"EA030003",
x"20030000",
x"08000604",
x"20030001",
x"08000609",
x"EA030003",
x"20030001",
x"08000609",
x"20030000",
x"E8800003",
x"44000806",
x"0800060D",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000611",
x"44810001",
x"44150802",
x"44210002",
x"44191803",
x"47431801",
x"44031803",
x"47031801",
x"44031803",
x"46E31801",
x"44030003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"08000624",
x"44200006",
x"C4260018",
x"44C01802",
x"200300B4",
x"C4610000",
x"44611802",
x"E7E302A0",
x"200300B0",
x"C4630000",
x"C4250014",
x"44A31802",
x"E7E3029C",
x"44C21802",
x"44610802",
x"E7E10298",
x"E7E20288",
x"E7F00284",
x"44000807",
x"E7E10280",
x"44A00807",
x"44200002",
x"E7E00294",
x"44C03007",
x"E7E60290",
x"44220002",
x"E7E0028C",
x"C7E1011C",
x"C7E002A0",
x"44200001",
x"E7E00128",
x"C7E10118",
x"C7E0029C",
x"44200001",
x"E7E00124",
x"C7E10114",
x"C7E00298",
x"44200001",
x"E7E00120",
x"40210024",
x"C00000C2",
x"C00000CF",
x"20210024",
x"C427001C",
x"44071002",
x"E8500003",
x"44400806",
x"08000653",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000679",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800066A",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000665",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"0800066A",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"08000679",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000674",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"08000679",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"0800069C",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800068D",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000688",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"0800068D",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"0800069C",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000697",
x"443D0800",
x"40210024",
x"C0000A77",
x"20210024",
x"0800069C",
x"443D0801",
x"40210024",
x"C0000A77",
x"20210024",
x"C4240010",
x"E8800006",
x"EA020003",
x"20030000",
x"080006A2",
x"20030001",
x"080006A7",
x"EA020003",
x"20030001",
x"080006A7",
x"20030000",
x"E8800003",
x"44000806",
x"080006AB",
x"47A00801",
x"EAC10003",
x"44200006",
x"080006AF",
x"44810001",
x"44150802",
x"44210002",
x"44191803",
x"47431801",
x"44031803",
x"47031801",
x"44031803",
x"46E31801",
x"44030003",
x"46200001",
x"44200003",
x"C42A000C",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"080006C3",
x"44200006",
x"44000007",
x"E7E00130",
x"E4220020",
x"40210028",
x"C00000CF",
x"20210028",
x"C427001C",
x"44071802",
x"C4220020",
x"46C21001",
x"E8500003",
x"44400806",
x"080006D1",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080006F7",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080006E8",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080006E3",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"080006E8",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"080006F7",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080006F2",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"080006F7",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"0800071A",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800070B",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000706",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800070B",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"0800071A",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000715",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800071A",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"C4240010",
x"E8800006",
x"EA020003",
x"20030000",
x"08000720",
x"20030001",
x"08000725",
x"EA020003",
x"20030001",
x"08000725",
x"20030000",
x"E8800003",
x"44000806",
x"08000729",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800072D",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"C42A000C",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44002807",
x"08000741",
x"44002806",
x"E8700003",
x"44600806",
x"08000745",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"0800076B",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800075C",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000757",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800075C",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"0800076B",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000766",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800076B",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"0800078E",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800077F",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800077A",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800077F",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"0800078E",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000789",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"0800078E",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"E8800006",
x"EA030003",
x"20030000",
x"08000793",
x"20030001",
x"08000798",
x"EA030003",
x"20030001",
x"08000798",
x"20030000",
x"E8800003",
x"44000806",
x"0800079C",
x"47A00801",
x"EAC10003",
x"44200006",
x"080007A0",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"080007B3",
x"44200006",
x"44A00002",
x"E7E00134",
x"46C31001",
x"E8500003",
x"44400806",
x"080007BA",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080007E0",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080007D1",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007CC",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"080007D1",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"080007E0",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007DB",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"080007E0",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"08000803",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080007F4",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007EF",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"080007F4",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"08000803",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007FE",
x"443D0800",
x"40210028",
x"C0000A77",
x"20210028",
x"08000803",
x"443D0801",
x"40210028",
x"C0000A77",
x"20210028",
x"E8800006",
x"EA020003",
x"20030000",
x"08000808",
x"20030001",
x"0800080D",
x"EA020003",
x"20030001",
x"0800080D",
x"20030000",
x"E8800003",
x"44000806",
x"08000811",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000815",
x"44810001",
x"44150002",
x"44001002",
x"44590803",
x"47410801",
x"44410803",
x"47010801",
x"44410803",
x"46E10801",
x"44410803",
x"46210801",
x"44010003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"08000828",
x"44200006",
x"44A00002",
x"E7E0012C",
x"40210028",
x"C00000CF",
x"E7E00138",
x"20080000",
x"C0000ED4",
x"20030000",
x"C000131B",
x"20040000",
x"C0001302",
x"AFE30204",
x"20030050",
x"04600001",
x"20030036",
x"04600001",
x"2003000A",
x"04600001",
x"8FE40258",
x"C0000BB4",
x"20030020",
x"04600001",
x"8FE40254",
x"C0000BB4",
x"20030020",
x"04600001",
x"200400FF",
x"C0000BB4",
x"2003000A",
x"04600001",
x"20060078",
x"20030003",
x"AFE2093C",
x"43E20904",
x"46000006",
x"C0000048",
x"20670000",
x"8FE2093C",
x"8FE3001C",
x"43E40904",
x"C000003F",
x"20640000",
x"AFE40908",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"20640000",
x"20C30000",
x"C000003F",
x"AFE302BC",
x"8FE602BC",
x"20030003",
x"AFE2093C",
x"43E20914",
x"46000006",
x"C0000048",
x"20670000",
x"8FE2093C",
x"8FE3001C",
x"43E40914",
x"C000003F",
x"20640000",
x"AFE40918",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE28",
x"20030003",
x"AFE2093C",
x"43E20924",
x"46000006",
x"C0000048",
x"20670000",
x"8FE2093C",
x"8FE3001C",
x"43E40924",
x"C000003F",
x"20640000",
x"AFE40928",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE2C",
x"20030003",
x"AFE2093C",
x"43E20934",
x"46000006",
x"C0000048",
x"20670000",
x"8FE2093C",
x"8FE3001C",
x"43E40934",
x"C000003F",
x"20640000",
x"AFE40938",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE30",
x"20070073",
x"C0003291",
x"20080003",
x"C00032EA",
x"20030009",
x"20080000",
x"200C0000",
x"C0000081",
x"20210028",
x"200300AC",
x"C4640000",
x"44040002",
x"200300A8",
x"C4630000",
x"44030001",
x"20030004",
x"E4200024",
x"4021002C",
x"C0000081",
x"2021002C",
x"44000806",
x"44240802",
x"44231001",
x"20040000",
x"C4200024",
x"E4230028",
x"E424002C",
x"E4210030",
x"21830000",
x"21050000",
x"46000806",
x"46002806",
x"40210038",
x"C0002FB7",
x"20210038",
x"200300A4",
x"C4650000",
x"C4210030",
x"44251000",
x"20040000",
x"20030002",
x"C4200024",
x"E4250034",
x"21050000",
x"46000806",
x"46002806",
x"4021003C",
x"C0002FB7",
x"2021003C",
x"20030003",
x"20050001",
x"AC250038",
x"40210040",
x"C0000081",
x"20210040",
x"44000806",
x"C424002C",
x"44240802",
x"C4230028",
x"44231001",
x"20040000",
x"C4200024",
x"8C250038",
x"E421003C",
x"21830000",
x"46000806",
x"46002806",
x"40210044",
x"C0002FB7",
x"20210044",
x"C4250034",
x"C421003C",
x"44251000",
x"20040000",
x"20080002",
x"C4200024",
x"8C250038",
x"21030000",
x"46000806",
x"46002806",
x"40210044",
x"C0002FB7",
x"20210044",
x"20030002",
x"20050002",
x"AC250040",
x"40210048",
x"C0000081",
x"20210048",
x"44000806",
x"C424002C",
x"44240802",
x"C4230028",
x"44231001",
x"20040000",
x"C4200024",
x"8C250040",
x"E4210044",
x"21830000",
x"46000806",
x"46002806",
x"4021004C",
x"C0002FB7",
x"2021004C",
x"C4250034",
x"C4210044",
x"44251000",
x"20040000",
x"C4200024",
x"8C250040",
x"21030000",
x"46000806",
x"46002806",
x"4021004C",
x"C0002FB7",
x"2021004C",
x"200A0001",
x"20090003",
x"C4200024",
x"21880000",
x"4021004C",
x"C00030B3",
x"200D0008",
x"200C0002",
x"20080004",
x"C000315E",
x"8FEB02BC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"200C0070",
x"C00033AD",
x"200D0003",
x"C000340E",
x"C7E00134",
x"E7E002DC",
x"C7E00130",
x"E7E002D8",
x"C7E0012C",
x"E7E002D4",
x"8FE3001C",
x"40650001",
x"43E702DC",
x"43E603CC",
x"C000132A",
x"2021004C",
x"8FE3001C",
x"40660001",
x"68C000D6",
x"A0C30002",
x"03E31820",
x"8C630110",
x"8C64FFF8",
x"20050002",
x"488500CF",
x"8C64FFE4",
x"C4800000",
x"E8110002",
x"08000A1E",
x"8C65FFFC",
x"48BC0084",
x"A0CB0002",
x"8FEC06B8",
x"C4800000",
x"46206001",
x"C7E10134",
x"44205807",
x"C7EA0130",
x"45405007",
x"C7E9012C",
x"45204807",
x"216E0001",
x"20030003",
x"46000006",
x"4021004C",
x"C0000048",
x"2021004C",
x"20640000",
x"8FE3001C",
x"AC240048",
x"40210050",
x"C000003F",
x"20210050",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240048",
x"ACA40000",
x"E4810000",
x"E48AFFFC",
x"E489FFF8",
x"8FE6001C",
x"40CD0001",
x"AC25004C",
x"21A50000",
x"20660000",
x"20870000",
x"40210054",
x"C000132A",
x"20210054",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C25004C",
x"AC65FFFC",
x"AC6E0000",
x"A1840002",
x"03E42020",
x"AC8306B4",
x"21920001",
x"216E0002",
x"C7E10130",
x"20030003",
x"46000006",
x"40210054",
x"C0000048",
x"20210054",
x"20640000",
x"8FE3001C",
x"AC240050",
x"40210058",
x"C000003F",
x"20210058",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240050",
x"ACA40000",
x"E48B0000",
x"E481FFFC",
x"E489FFF8",
x"8FE6001C",
x"40CD0001",
x"AC250054",
x"21A50000",
x"20660000",
x"20870000",
x"4021005C",
x"C000132A",
x"2021005C",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C250054",
x"AC65FFFC",
x"AC6E0000",
x"A2440002",
x"03E42020",
x"AC8306B4",
x"218E0002",
x"216D0003",
x"C7E1012C",
x"20030003",
x"46000006",
x"4021005C",
x"C0000048",
x"2021005C",
x"20640000",
x"8FE3001C",
x"AC240058",
x"40210060",
x"C000003F",
x"20210060",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240058",
x"ACA40000",
x"E48B0000",
x"E48AFFFC",
x"E481FFF8",
x"8FE6001C",
x"40CB0001",
x"AC25005C",
x"21650000",
x"20660000",
x"20870000",
x"40210064",
x"C000132A",
x"20210064",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C25005C",
x"AC65FFFC",
x"AC6D0000",
x"A1C40002",
x"03E42020",
x"AC8306B4",
x"21830003",
x"AFE306B8",
x"08000A1E",
x"20040002",
x"48A40043",
x"A0C40002",
x"208C0001",
x"8FED06B8",
x"46204801",
x"8C63FFF0",
x"C7E70134",
x"C4650000",
x"44E51002",
x"C7E10130",
x"C466FFFC",
x"44260002",
x"44402000",
x"C7E2012C",
x"C460FFF8",
x"44401802",
x"44831800",
x"C42A000C",
x"45452002",
x"44832002",
x"44872801",
x"45462002",
x"44832002",
x"44812001",
x"45400002",
x"44030002",
x"44020801",
x"20030003",
x"46000006",
x"40210064",
x"C0000048",
x"20210064",
x"20640000",
x"8FE3001C",
x"AC240060",
x"40210068",
x"C000003F",
x"20210068",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240060",
x"ACA40000",
x"E4850000",
x"E484FFFC",
x"E481FFF8",
x"8FE6001C",
x"40CB0001",
x"AC250064",
x"21650000",
x"20660000",
x"20870000",
x"4021006C",
x"C000132A",
x"2021006C",
x"20430000",
x"2042000C",
x"E469FFF8",
x"8C250064",
x"AC65FFFC",
x"AC6C0000",
x"A1A40002",
x"03E42020",
x"AC8306B4",
x"21A30001",
x"AFE306B8",
x"08000A1E",
x"08000A1F",
x"08000A20",
x"20080000",
x"C7E30264",
x"8FE3025C",
x"00031822",
x"4021006C",
x"C0000081",
x"2021006C",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"8C300008",
x"22070000",
x"4021006C",
x"C0002DD9",
x"2021006C",
x"200A0000",
x"20080002",
x"8FE30254",
x"69430002",
x"08000A75",
x"40630001",
x"AC2A0068",
x"69430002",
x"08000A5F",
x"20040001",
x"C7E30264",
x"8FE3025C",
x"00831822",
x"40210070",
x"C0000081",
x"20210070",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"8C2F0004",
x"21E70000",
x"40210070",
x"C0002DD9",
x"20210070",
x"20060000",
x"8C2A0068",
x"8C310000",
x"8C300008",
x"8C2F0004",
x"21E80000",
x"22070000",
x"22290000",
x"40210070",
x"C0002E50",
x"20210070",
x"200A0001",
x"20030004",
x"8C300008",
x"8C2F0004",
x"8C310000",
x"22280000",
x"21E90000",
x"22070000",
x"40210070",
x"C0002EBB",
x"20210070",
x"20000000",
x"0000003F",
x"EBA10037",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1001B",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA1001B",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000A77",
x"443D0801",
x"08000A77",
x"012A1820",
x"A8650001",
x"00A63818",
x"01491822",
x"6B830003",
x"21230000",
x"E0000000",
x"68E40068",
x"48E40003",
x"20A30000",
x"E0000000",
x"01251820",
x"A8670001",
x"00E64018",
x"00A91822",
x"6B830003",
x"21230000",
x"E0000000",
x"69040030",
x"49040003",
x"20E30000",
x"E0000000",
x"01271820",
x"A8680001",
x"01062818",
x"00E91822",
x"6B830003",
x"21230000",
x"E0000000",
x"68A40014",
x"48A40003",
x"21030000",
x"E0000000",
x"01281820",
x"A8650001",
x"00A63818",
x"01091822",
x"6B830003",
x"21230000",
x"E0000000",
x"68E40006",
x"48E40003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"08000AE1",
x"210A0000",
x"20A90000",
x"08000AE1",
x"01071820",
x"A8650001",
x"00A64818",
x"00E81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"21090000",
x"08000AE1",
x"20EA0000",
x"20A90000",
x"08000AE1",
x"00E51820",
x"A8680001",
x"01064818",
x"00A71822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240015",
x"49240003",
x"21030000",
x"E0000000",
x"00E81820",
x"A8650001",
x"00A64818",
x"01071822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000AE1",
x"210A0000",
x"20A90000",
x"08000AE1",
x"01051820",
x"A8670001",
x"00E64818",
x"00A81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20E30000",
x"E0000000",
x"20EA0000",
x"21090000",
x"08000AE1",
x"20AA0000",
x"20E90000",
x"08000AE1",
x"00AA1820",
x"A8680001",
x"01063818",
x"01451822",
x"6B830003",
x"20A30000",
x"E0000000",
x"68E40031",
x"48E40003",
x"21030000",
x"E0000000",
x"00A81820",
x"A8670001",
x"00E64818",
x"01051822",
x"6B830003",
x"20A30000",
x"E0000000",
x"69240015",
x"49240003",
x"20E30000",
x"E0000000",
x"00A71820",
x"A8680001",
x"01064818",
x"00E51822",
x"6B830003",
x"20A30000",
x"E0000000",
x"69240007",
x"49240003",
x"21030000",
x"E0000000",
x"210A0000",
x"20A90000",
x"08000AE1",
x"20EA0000",
x"21090000",
x"08000AE1",
x"00E81820",
x"A8650001",
x"00A64818",
x"01071822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000AE1",
x"210A0000",
x"20A90000",
x"08000AE1",
x"010A1820",
x"A8670001",
x"00E62818",
x"01481822",
x"6B830003",
x"21030000",
x"E0000000",
x"68A40015",
x"48A40003",
x"20E30000",
x"E0000000",
x"01071820",
x"A8650001",
x"00A64818",
x"00E81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"21090000",
x"08000AE1",
x"20EA0000",
x"20A90000",
x"08000AE1",
x"00EA1820",
x"A8650001",
x"00A64018",
x"01471822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69040007",
x"49040003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000AE1",
x"20A90000",
x"08000AE1",
x"6880031C",
x"3C6005F5",
x"1C60E100",
x"68640006",
x"48640003",
x"20050001",
x"08000BBC",
x"20050000",
x"08000BC6",
x"3C600BEB",
x"1C60C200",
x"68640006",
x"48640003",
x"20050002",
x"08000BC4",
x"20050001",
x"08000BC6",
x"20050002",
x"3C6005F5",
x"1C60E100",
x"00A31818",
x"00832022",
x"68050003",
x"200D0000",
x"08000BD1",
x"20030030",
x"00651820",
x"04600001",
x"200D0001",
x"3CC00098",
x"1CC09680",
x"200C0000",
x"200A000A",
x"20090005",
x"3CA002FA",
x"1CA0F080",
x"AC240000",
x"68A40030",
x"48A40003",
x"20030005",
x"08000C08",
x"200B0002",
x"3CA00131",
x"1CA02D00",
x"68A40016",
x"48A40003",
x"20030002",
x"08000BF5",
x"20090001",
x"3CA00098",
x"1CA09680",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000BF0",
x"212A0000",
x"21890000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000BF5",
x"216A0000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C08",
x"200A0003",
x"3CA001C9",
x"1CA0C380",
x"68A40009",
x"48A40003",
x"20030003",
x"08000C01",
x"21690000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C08",
x"215B0000",
x"212A0000",
x"23690000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C31",
x"200B0007",
x"3CA0042C",
x"1CA01D80",
x"68A40015",
x"48A40003",
x"20030007",
x"08000C20",
x"200A0006",
x"3CA00393",
x"1CA08700",
x"68A40008",
x"48A40003",
x"20030006",
x"08000C1A",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C20",
x"21490000",
x"216A0000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C31",
x"20090008",
x"3CA004C4",
x"1CA0B400",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000C2D",
x"212A0000",
x"21690000",
x"40210008",
x"C0000AE1",
x"20210008",
x"08000C31",
x"40210008",
x"C0000AE1",
x"20210008",
x"3CA00098",
x"1CA09680",
x"00652818",
x"8C240000",
x"00852022",
x"68030009",
x"49A00003",
x"200E0000",
x"08000C3E",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"08000C43",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"3CC0000F",
x"1CC04240",
x"200C0000",
x"200A000A",
x"20090005",
x"3CA0004C",
x"1CA04B40",
x"AC240004",
x"68A40030",
x"48A40003",
x"20030005",
x"08000C7A",
x"200B0002",
x"3CA0001E",
x"1CA08480",
x"68A40016",
x"48A40003",
x"20030002",
x"08000C67",
x"20090001",
x"3CA0000F",
x"1CA04240",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000C62",
x"212A0000",
x"21890000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000C67",
x"216A0000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000C7A",
x"200A0003",
x"3CA0002D",
x"1CA0C6C0",
x"68A40009",
x"48A40003",
x"20030003",
x"08000C73",
x"21690000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000C7A",
x"215B0000",
x"212A0000",
x"23690000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000CA3",
x"200B0007",
x"3CA0006A",
x"1CA0CFC0",
x"68A40015",
x"48A40003",
x"20030007",
x"08000C92",
x"200A0006",
x"3CA0005B",
x"1CA08D80",
x"68A40008",
x"48A40003",
x"20030006",
x"08000C8C",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000C92",
x"21490000",
x"216A0000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000CA3",
x"20090008",
x"3CA0007A",
x"1CA01200",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000C9F",
x"212A0000",
x"21690000",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"08000CA3",
x"4021000C",
x"C0000AE1",
x"2021000C",
x"3CA0000F",
x"1CA04240",
x"00652818",
x"8C240004",
x"00852022",
x"68030009",
x"49C00003",
x"200D0000",
x"08000CB0",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"08000CB5",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"3CC00001",
x"1CC086A0",
x"200C0000",
x"200A000A",
x"20090005",
x"3CA00007",
x"1CA0A120",
x"AC240008",
x"68A40030",
x"48A40003",
x"20030005",
x"08000CEC",
x"200B0002",
x"3CA00003",
x"1CA00D40",
x"68A40016",
x"48A40003",
x"20030002",
x"08000CD9",
x"20090001",
x"3CA00001",
x"1CA086A0",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000CD4",
x"212A0000",
x"21890000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000CD9",
x"216A0000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000CEC",
x"200A0003",
x"3CA00004",
x"1CA093E0",
x"68A40009",
x"48A40003",
x"20030003",
x"08000CE5",
x"21690000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000CEC",
x"215B0000",
x"212A0000",
x"23690000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000D15",
x"200B0007",
x"3CA0000A",
x"1CA0AE60",
x"68A40015",
x"48A40003",
x"20030007",
x"08000D04",
x"200A0006",
x"3CA00009",
x"1CA027C0",
x"68A40008",
x"48A40003",
x"20030006",
x"08000CFE",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000D04",
x"21490000",
x"216A0000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000D15",
x"20090008",
x"3CA0000C",
x"1CA03500",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000D11",
x"212A0000",
x"21690000",
x"40210010",
x"C0000AE1",
x"20210010",
x"08000D15",
x"40210010",
x"C0000AE1",
x"20210010",
x"3CA00001",
x"1CA086A0",
x"00652818",
x"8C240008",
x"00852022",
x"68030009",
x"49A00003",
x"200E0000",
x"08000D22",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"08000D27",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"20062710",
x"200C0000",
x"200A000A",
x"20090005",
x"3CA00000",
x"1CA0C350",
x"AC24000C",
x"68A4002D",
x"48A40003",
x"20030005",
x"08000D5A",
x"200B0002",
x"20054E20",
x"68A40015",
x"48A40003",
x"20030002",
x"08000D48",
x"20090001",
x"20052710",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000D43",
x"212A0000",
x"21890000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D48",
x"216A0000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D5A",
x"200A0003",
x"20057530",
x"68A40009",
x"48A40003",
x"20030003",
x"08000D53",
x"21690000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D5A",
x"215B0000",
x"212A0000",
x"23690000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D83",
x"200B0007",
x"3CA00001",
x"1CA01170",
x"68A40015",
x"48A40003",
x"20030007",
x"08000D72",
x"200A0006",
x"3CA00000",
x"1CA0EA60",
x"68A40008",
x"48A40003",
x"20030006",
x"08000D6C",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D72",
x"21490000",
x"216A0000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D83",
x"20090008",
x"3CA00001",
x"1CA03880",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000D7F",
x"212A0000",
x"21690000",
x"40210014",
x"C0000AE1",
x"20210014",
x"08000D83",
x"40210014",
x"C0000AE1",
x"20210014",
x"20052710",
x"00652818",
x"8C24000C",
x"00852022",
x"68030009",
x"49C00003",
x"200D0000",
x"08000D8F",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"08000D94",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"200603E8",
x"200C0000",
x"200A000A",
x"20090005",
x"20051388",
x"AC240010",
x"68A4002D",
x"48A40003",
x"20030005",
x"08000DC6",
x"200B0002",
x"200507D0",
x"68A40015",
x"48A40003",
x"20030002",
x"08000DB4",
x"20090001",
x"200503E8",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000DAF",
x"212A0000",
x"21890000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DB4",
x"216A0000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DC6",
x"200A0003",
x"20050BB8",
x"68A40009",
x"48A40003",
x"20030003",
x"08000DBF",
x"21690000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DC6",
x"215B0000",
x"212A0000",
x"23690000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DEC",
x"200B0007",
x"20051B58",
x"68A40014",
x"48A40003",
x"20030007",
x"08000DDC",
x"200A0006",
x"20051770",
x"68A40008",
x"48A40003",
x"20030006",
x"08000DD6",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DDC",
x"21490000",
x"216A0000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DEC",
x"20090008",
x"20051F40",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000DE8",
x"212A0000",
x"21690000",
x"40210018",
x"C0000AE1",
x"20210018",
x"08000DEC",
x"40210018",
x"C0000AE1",
x"20210018",
x"606503E8",
x"8C240010",
x"00852022",
x"68030009",
x"49A00003",
x"200E0000",
x"08000DF7",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"08000DFC",
x"20050030",
x"00A31820",
x"04600001",
x"200E0001",
x"20060064",
x"200C0000",
x"200A000A",
x"20090005",
x"200501F4",
x"AC240014",
x"68A4002D",
x"48A40003",
x"20030005",
x"08000E2E",
x"200B0002",
x"200500C8",
x"68A40015",
x"48A40003",
x"20030002",
x"08000E1C",
x"20090001",
x"20050064",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000E17",
x"212A0000",
x"21890000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E1C",
x"216A0000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E2E",
x"200A0003",
x"2005012C",
x"68A40009",
x"48A40003",
x"20030003",
x"08000E27",
x"21690000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E2E",
x"215B0000",
x"212A0000",
x"23690000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E54",
x"200B0007",
x"200502BC",
x"68A40014",
x"48A40003",
x"20030007",
x"08000E44",
x"200A0006",
x"20050258",
x"68A40008",
x"48A40003",
x"20030006",
x"08000E3E",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E44",
x"21490000",
x"216A0000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E54",
x"20090008",
x"20050320",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000E50",
x"212A0000",
x"21690000",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"08000E54",
x"4021001C",
x"C0000AE1",
x"2021001C",
x"60650064",
x"8C240014",
x"00852022",
x"68030009",
x"49C00003",
x"200D0000",
x"08000E5F",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"08000E64",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"2006000A",
x"200C0000",
x"200A000A",
x"20090005",
x"20050032",
x"AC240018",
x"68A4002D",
x"48A40003",
x"20030005",
x"08000E96",
x"200B0002",
x"20050014",
x"68A40015",
x"48A40003",
x"20030002",
x"08000E84",
x"20090001",
x"2005000A",
x"68A4000A",
x"48A40003",
x"20030001",
x"08000E7F",
x"212A0000",
x"21890000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000E84",
x"216A0000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000E96",
x"200A0003",
x"2005001E",
x"68A40009",
x"48A40003",
x"20030003",
x"08000E8F",
x"21690000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000E96",
x"215B0000",
x"212A0000",
x"23690000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000EBC",
x"200B0007",
x"20050046",
x"68A40014",
x"48A40003",
x"20030007",
x"08000EAC",
x"200A0006",
x"2005003C",
x"68A40008",
x"48A40003",
x"20030006",
x"08000EA6",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000EAC",
x"21490000",
x"216A0000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000EBC",
x"20090008",
x"20050050",
x"68A4000A",
x"48A40003",
x"20030008",
x"08000EB8",
x"212A0000",
x"21690000",
x"40210020",
x"C0000AE1",
x"20210020",
x"08000EBC",
x"40210020",
x"C0000AE1",
x"20210020",
x"6065000A",
x"8C240018",
x"00852022",
x"68030009",
x"49A00003",
x"20050000",
x"08000EC7",
x"20050030",
x"00A31820",
x"04600001",
x"20050001",
x"08000ECC",
x"20050030",
x"00A31820",
x"04600001",
x"20050001",
x"20030030",
x"00641820",
x"04600001",
x"E0000000",
x"2003002D",
x"04600001",
x"00042022",
x"08000BB4",
x"2003003C",
x"69030002",
x"E0000000",
x"AC280000",
x"40210008",
x"C00000C2",
x"20210008",
x"206B0000",
x"497D0003",
x"20030000",
x"080012E5",
x"AC2B0004",
x"4021000C",
x"C00000C2",
x"2021000C",
x"20660000",
x"AC260008",
x"40210010",
x"C00000C2",
x"20210010",
x"206C0000",
x"AC2C000C",
x"40210014",
x"C00000C2",
x"20670000",
x"20030003",
x"46000006",
x"C0000048",
x"20210014",
x"20650000",
x"AC270010",
x"AC250014",
x"4021001C",
x"C00000CF",
x"2021001C",
x"8C250014",
x"E4A00000",
x"4021001C",
x"C00000CF",
x"2021001C",
x"8C250014",
x"E4A0FFFC",
x"4021001C",
x"C00000CF",
x"2021001C",
x"8C250014",
x"E4A0FFF8",
x"20030003",
x"46000006",
x"4021001C",
x"C0000048",
x"2021001C",
x"206A0000",
x"AC2A0018",
x"40210020",
x"C00000CF",
x"20210020",
x"8C2A0018",
x"E5400000",
x"40210020",
x"C00000CF",
x"20210020",
x"8C2A0018",
x"E540FFFC",
x"40210020",
x"C00000CF",
x"20210020",
x"8C2A0018",
x"E540FFF8",
x"40210020",
x"C00000CF",
x"44001006",
x"20030002",
x"46000006",
x"C0000048",
x"20210020",
x"206D0000",
x"E422001C",
x"AC2D0020",
x"40210028",
x"C00000CF",
x"20210028",
x"8C2D0020",
x"E5A00000",
x"40210028",
x"C00000CF",
x"20210028",
x"8C2D0020",
x"E5A0FFFC",
x"20030003",
x"46000006",
x"40210028",
x"C0000048",
x"20210028",
x"206E0000",
x"AC2E0024",
x"4021002C",
x"C00000CF",
x"2021002C",
x"8C2E0024",
x"E5C00000",
x"4021002C",
x"C00000CF",
x"2021002C",
x"8C2E0024",
x"E5C0FFFC",
x"4021002C",
x"C00000CF",
x"2021002C",
x"8C2E0024",
x"E5C0FFF8",
x"20030003",
x"46000006",
x"4021002C",
x"C0000048",
x"2021002C",
x"8C270010",
x"48E00002",
x"08000F63",
x"AC230028",
x"40210030",
x"C00000CF",
x"20210030",
x"200400CC",
x"C4810000",
x"44010002",
x"8C230028",
x"E4600000",
x"E421002C",
x"40210034",
x"C00000CF",
x"20210034",
x"C421002C",
x"44010002",
x"8C230028",
x"E460FFFC",
x"40210034",
x"C00000CF",
x"20210034",
x"C421002C",
x"44010002",
x"8C230028",
x"E460FFF8",
x"200F0002",
x"8C260008",
x"48CF0003",
x"200F0001",
x"08000F6D",
x"C422001C",
x"E8500003",
x"200F0000",
x"08000F6D",
x"200F0001",
x"20090004",
x"AC230028",
x"21230000",
x"46000006",
x"40210034",
x"C0000048",
x"20210034",
x"20690000",
x"20440000",
x"2042002C",
x"AC89FFD8",
x"8C230028",
x"AC83FFDC",
x"8C2E0024",
x"AC8EFFE0",
x"8C2D0020",
x"AC8DFFE4",
x"AC8FFFE8",
x"8C2A0018",
x"AC8AFFEC",
x"8C250014",
x"AC85FFF0",
x"8C270010",
x"AC87FFF4",
x"8C2C000C",
x"AC8CFFF8",
x"AC86FFFC",
x"8C2B0004",
x"AC8B0000",
x"8C280000",
x"A1090002",
x"03E94820",
x"AD240110",
x"20040003",
x"48C40032",
x"C4A10000",
x"C830000D",
x"C8300008",
x"EA010004",
x"200400A0",
x"C4800000",
x"08000F99",
x"200400C8",
x"C4800000",
x"08000F9B",
x"46000006",
x"44210802",
x"44010003",
x"08000F9F",
x"46000006",
x"E4A00000",
x"C4A1FFFC",
x"C830000D",
x"C8300008",
x"EA010004",
x"200400A0",
x"C4800000",
x"08000FA9",
x"200400C8",
x"C4800000",
x"08000FAB",
x"46000006",
x"44210802",
x"44010003",
x"08000FAF",
x"46000006",
x"E4A0FFFC",
x"C4A1FFF8",
x"C830000D",
x"C8300008",
x"EA010004",
x"200400A0",
x"C4800000",
x"08000FB9",
x"200400C8",
x"C4800000",
x"08000FBB",
x"46000006",
x"44210802",
x"44010003",
x"08000FBF",
x"46000006",
x"E4A0FFF8",
x"08000FDE",
x"20040002",
x"48C4001C",
x"C4A10000",
x"44211802",
x"C4A0FFFC",
x"44000002",
x"44601800",
x"C4A0FFF8",
x"44000002",
x"44600000",
x"44001804",
x"C8700007",
x"C422001C",
x"E8500003",
x"46830003",
x"08000FD2",
x"46230003",
x"08000FD5",
x"200400C8",
x"C4800000",
x"44200802",
x"E4A10000",
x"C4A1FFFC",
x"44200802",
x"E4A1FFFC",
x"C4A1FFF8",
x"44200002",
x"E4A0FFF8",
x"08000FDE",
x"48E00002",
x"080012E4",
x"C4630000",
x"46C31001",
x"200400F0",
x"C4840000",
x"200400EC",
x"C48E0000",
x"E8500003",
x"44400806",
x"08000FEA",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001010",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001001",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000FFC",
x"443D0800",
x"40210034",
x"C0000A77",
x"20210034",
x"08001001",
x"443D0801",
x"40210034",
x"C0000A77",
x"20210034",
x"08001010",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800100B",
x"443D0800",
x"40210034",
x"C0000A77",
x"20210034",
x"08001010",
x"443D0801",
x"40210034",
x"C0000A77",
x"20210034",
x"08001033",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001024",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800101F",
x"443D0800",
x"40210034",
x"C0000A77",
x"20210034",
x"08001024",
x"443D0801",
x"40210034",
x"C0000A77",
x"20210034",
x"08001033",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800102E",
x"443D0800",
x"40210034",
x"C0000A77",
x"20210034",
x"08001033",
x"443D0801",
x"40210034",
x"C0000A77",
x"20210034",
x"E8800006",
x"EA020003",
x"20040000",
x"08001038",
x"20040001",
x"0800103D",
x"EA020003",
x"20040001",
x"0800103D",
x"20040000",
x"E8800003",
x"44000806",
x"08001041",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001045",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48800003",
x"44007807",
x"08001058",
x"44007806",
x"E8700003",
x"44600806",
x"0800105C",
x"44600807",
x"E42F0030",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001083",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001074",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800106F",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001074",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001083",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800107E",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001083",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"080010A6",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001097",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001092",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001097",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"080010A6",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080010A1",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080010A6",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"E8800006",
x"EA030003",
x"20040000",
x"080010AB",
x"20040001",
x"080010B0",
x"EA030003",
x"20040001",
x"080010B0",
x"20040000",
x"E8800003",
x"44000806",
x"080010B4",
x"47A00801",
x"EAC10003",
x"44200006",
x"080010B8",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48800003",
x"44003807",
x"080010CB",
x"44003806",
x"C463FFFC",
x"46C31001",
x"E8500003",
x"44400806",
x"080010D1",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080010F7",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080010E8",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080010E3",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080010E8",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"080010F7",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080010F2",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080010F7",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"0800111A",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800110B",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001106",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800110B",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"0800111A",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001115",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800111A",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"E8800006",
x"EA020003",
x"20040000",
x"0800111F",
x"20040001",
x"08001124",
x"EA020003",
x"20040001",
x"08001124",
x"20040000",
x"E8800003",
x"44000806",
x"08001128",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800112C",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200803",
x"45C10002",
x"44210802",
x"46210800",
x"44010003",
x"48800003",
x"44006807",
x"0800113F",
x"44006806",
x"E8700003",
x"44600806",
x"08001143",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001169",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800115A",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001155",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800115A",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001169",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001164",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001169",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"0800118C",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800117D",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001178",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800117D",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"0800118C",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001187",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800118C",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"E8800006",
x"EA030003",
x"20040000",
x"08001191",
x"20040001",
x"08001196",
x"EA030003",
x"20040001",
x"08001196",
x"20040000",
x"E8800003",
x"44000806",
x"0800119A",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800119E",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200803",
x"45C10002",
x"44210802",
x"46210800",
x"44010003",
x"48800003",
x"44004807",
x"080011B1",
x"44004806",
x"C463FFF8",
x"46C31001",
x"E8500003",
x"44400806",
x"080011B7",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080011DD",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080011CE",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080011C9",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080011CE",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"080011DD",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080011D8",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080011DD",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001200",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080011F1",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080011EC",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"080011F1",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001200",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080011FB",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001200",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"E8800006",
x"EA020003",
x"20040000",
x"08001205",
x"20040001",
x"0800120A",
x"EA020003",
x"20040001",
x"0800120A",
x"20040000",
x"E8800003",
x"44000806",
x"0800120E",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001212",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48800003",
x"44001007",
x"08001225",
x"44001006",
x"E8700003",
x"44600806",
x"08001229",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"0800124F",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001240",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800123B",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001240",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"0800124F",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800124A",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"0800124F",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001272",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001263",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800125E",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001263",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"08001272",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800126D",
x"443D0800",
x"40210038",
x"C0000A77",
x"20210038",
x"08001272",
x"443D0801",
x"40210038",
x"C0000A77",
x"20210038",
x"E8800006",
x"EA030003",
x"20040000",
x"08001277",
x"20040001",
x"0800127C",
x"EA030003",
x"20040001",
x"0800127C",
x"20040000",
x"E8800003",
x"44000806",
x"08001280",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001284",
x"44810001",
x"44150802",
x"44210002",
x"44191803",
x"47431801",
x"44031803",
x"47031801",
x"44031803",
x"46E31801",
x"44030003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200803",
x"48800003",
x"44200007",
x"08001297",
x"44200006",
x"45A26002",
x"44E92802",
x"44A21802",
x"C42F0030",
x"45E00802",
x"44615001",
x"45E90802",
x"44222002",
x"44E01802",
x"44833000",
x"45A05802",
x"44A02002",
x"45E21802",
x"44834000",
x"44200802",
x"44E20002",
x"44202801",
x"45204807",
x"44ED3802",
x"45ED2002",
x"C4A00000",
x"C4A2FFFC",
x"C4A3FFF8",
x"458C0802",
x"44016802",
x"456B0802",
x"44410802",
x"45A16800",
x"45290802",
x"44610802",
x"45A10800",
x"E4A10000",
x"454A0802",
x"44016802",
x"45080802",
x"44410802",
x"45A16800",
x"44E70802",
x"44610802",
x"45A10800",
x"E4A1FFFC",
x"44C60802",
x"44016802",
x"44A50802",
x"44410802",
x"45A16800",
x"44840802",
x"44610802",
x"45A10800",
x"E4A1FFF8",
x"440A0802",
x"44266802",
x"44480802",
x"44250802",
x"45A16800",
x"44670802",
x"44240802",
x"45A10800",
x"45C10802",
x"E4610000",
x"440C0802",
x"44263002",
x"444B0002",
x"44051002",
x"44C22800",
x"44691802",
x"44641002",
x"44A21000",
x"45C21002",
x"E462FFFC",
x"442A0802",
x"44080002",
x"44200800",
x"44670002",
x"44200000",
x"45C00002",
x"E460FFF8",
x"20030001",
x"48600004",
x"8C280000",
x"AFE8001C",
x"E0000000",
x"8C280000",
x"21080001",
x"08000ED4",
x"AC240000",
x"40210008",
x"C00000C2",
x"20210008",
x"20650000",
x"48BD0005",
x"8C240000",
x"20830001",
x"2004FFFF",
x"0800003F",
x"8C240000",
x"20830001",
x"AC250004",
x"20640000",
x"4021000C",
x"C00012EC",
x"2021000C",
x"8C240000",
x"A0840002",
x"8C250004",
x"6C642800",
x"E0000000",
x"20030000",
x"AC240000",
x"20640000",
x"40210008",
x"C00012EC",
x"20210008",
x"20660000",
x"8CC30000",
x"487D0005",
x"8C240000",
x"20830001",
x"20C40000",
x"0800003F",
x"8C240000",
x"20830001",
x"AC260004",
x"20640000",
x"4021000C",
x"C0001302",
x"2021000C",
x"8C240000",
x"A0840002",
x"8C260004",
x"6C643000",
x"E0000000",
x"20040000",
x"AC230000",
x"40210008",
x"C00012EC",
x"20210008",
x"20640000",
x"8C850000",
x"48BD0002",
x"E0000000",
x"8C230000",
x"A0650002",
x"03E52820",
x"ACA40200",
x"20630001",
x"0800131B",
x"68A000C6",
x"A0A30002",
x"03E31820",
x"8C690110",
x"8D23FFFC",
x"487C0042",
x"20030006",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E00000",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"0800133C",
x"200A0001",
x"8D28FFF0",
x"C5010000",
x"488A0003",
x"44200007",
x"08001342",
x"44200006",
x"E4600000",
x"C4E00000",
x"46200003",
x"E460FFFC",
x"08001348",
x"E470FFFC",
x"C4E0FFFC",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"0800134F",
x"200A0001",
x"8D28FFF0",
x"C501FFFC",
x"488A0003",
x"44200007",
x"08001355",
x"44200006",
x"E460FFF8",
x"C4E0FFFC",
x"46200003",
x"E460FFF4",
x"0800135B",
x"E470FFF4",
x"C4E0FFF8",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"08001362",
x"200A0001",
x"8D28FFF0",
x"C501FFF8",
x"488A0003",
x"44200007",
x"08001368",
x"44200006",
x"E460FFF0",
x"C4E0FFF8",
x"46200003",
x"E460FFEC",
x"0800136E",
x"E470FFEC",
x"A0A40002",
x"6CC41800",
x"080013EE",
x"20040002",
x"48640026",
x"20030004",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E10000",
x"8D24FFF0",
x"C4800000",
x"44201002",
x"C4E1FFFC",
x"C480FFFC",
x"44200002",
x"44401000",
x"C4E1FFF8",
x"C480FFF8",
x"44200002",
x"44400000",
x"EA000003",
x"E4700000",
x"08001395",
x"46800803",
x"E4610000",
x"C4810000",
x"44200803",
x"44200807",
x"E461FFFC",
x"C481FFFC",
x"44200803",
x"44200807",
x"E461FFF8",
x"C481FFF8",
x"44200003",
x"44000007",
x"E460FFF4",
x"A0A40002",
x"6CC41800",
x"080013EE",
x"20030005",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E00000",
x"C4E1FFFC",
x"C4E2FFF8",
x"44001802",
x"8D24FFF0",
x"C4850000",
x"44652002",
x"44211802",
x"C486FFFC",
x"44661802",
x"44833800",
x"44421802",
x"C484FFF8",
x"44641802",
x"44E33800",
x"8D28FFF4",
x"49000003",
x"44E01806",
x"080013BD",
x"44224002",
x"8D24FFDC",
x"C4830000",
x"45031802",
x"44E34000",
x"44403802",
x"C483FFFC",
x"44E31802",
x"45034000",
x"44013802",
x"C483FFF8",
x"44E31802",
x"45031800",
x"44050002",
x"44000007",
x"44260802",
x"44200807",
x"44441002",
x"44401007",
x"E4630000",
x"49000005",
x"E460FFFC",
x"E461FFF8",
x"E462FFF4",
x"080013E8",
x"C4E5FFF8",
x"8D24FFDC",
x"C484FFFC",
x"44A43002",
x"C4E5FFFC",
x"C484FFF8",
x"44A42002",
x"44C42000",
x"44952002",
x"44040001",
x"E460FFFC",
x"C4E4FFF8",
x"C4800000",
x"44802802",
x"C4E40000",
x"C480FFF8",
x"44800002",
x"44A00000",
x"44150002",
x"44200001",
x"E460FFF8",
x"C4E1FFFC",
x"C4800000",
x"44202002",
x"C4E10000",
x"C480FFFC",
x"44200002",
x"44800000",
x"44150002",
x"44400001",
x"E460FFF4",
x"C8700004",
x"46230003",
x"E460FFF0",
x"080013EC",
x"A0A40002",
x"6CC41800",
x"40A50001",
x"0800132A",
x"E0000000",
x"6880009C",
x"A0850002",
x"03E52820",
x"8CA50110",
x"8CA8FFD8",
x"8CA7FFFC",
x"C4610000",
x"8CA6FFEC",
x"C4C00000",
x"44200001",
x"E5000000",
x"C461FFFC",
x"C4C0FFFC",
x"44200001",
x"E500FFFC",
x"C461FFF8",
x"C4C0FFF8",
x"44200001",
x"E500FFF8",
x"20060002",
x"48E6000F",
x"8CA5FFF0",
x"C5010000",
x"C503FFFC",
x"C502FFF8",
x"C4A00000",
x"44010802",
x"C4A0FFFC",
x"44030002",
x"44200800",
x"C4A0FFF8",
x"44020002",
x"44200000",
x"E500FFF4",
x"0800143D",
x"20060002",
x"68C70002",
x"0800143D",
x"C5020000",
x"C501FFFC",
x"C500FFF8",
x"44422002",
x"8CA6FFF0",
x"C4C30000",
x"44832802",
x"44212002",
x"C4C3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4C3FFF8",
x"44831802",
x"44A32000",
x"8CA6FFF4",
x"48C00003",
x"44801806",
x"08001437",
x"44202802",
x"8CA5FFDC",
x"C4A30000",
x"44A31802",
x"44832000",
x"44021802",
x"C4A0FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C4A0FFF8",
x"44201802",
x"44831800",
x"20050003",
x"48E50003",
x"44710001",
x"0800143C",
x"44600006",
x"E500FFF4",
x"40880001",
x"6900004E",
x"A1040002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C4610000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C461FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C461FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"0800148A",
x"20050002",
x"68A60002",
x"0800148A",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08001484",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08001489",
x"44600006",
x"E4E0FFF4",
x"41040001",
x"080013F1",
x"E0000000",
x"E0000000",
x"A0A30002",
x"4C833000",
x"48DD0003",
x"20030001",
x"E0000000",
x"A0C30002",
x"03E31820",
x"8C670110",
x"8CE3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CE6FFFC",
x"48DC0024",
x"E8100003",
x"44003006",
x"080014A3",
x"44003007",
x"8CE3FFF0",
x"C4600000",
x"E8C00003",
x"20060000",
x"080014B9",
x"E8500003",
x"44400006",
x"080014AC",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20060000",
x"080014B9",
x"E8300003",
x"44200006",
x"080014B4",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20060000",
x"080014B9",
x"20060001",
x"48C00007",
x"8CE3FFE8",
x"48600003",
x"20030001",
x"080014BF",
x"20030000",
x"080014C1",
x"8CE3FFE8",
x"08001502",
x"20030002",
x"48C30014",
x"8CE3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CE3FFE8",
x"E8100003",
x"20060000",
x"080014D2",
x"20060001",
x"48660003",
x"20030001",
x"080014D6",
x"20030000",
x"08001502",
x"44003802",
x"8CE3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CE3FFF4",
x"48600003",
x"44E03006",
x"080014F4",
x"44414002",
x"8CE3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48C30003",
x"44D10001",
x"080014F9",
x"44C00006",
x"8CE3FFE8",
x"E8100003",
x"20060000",
x"080014FE",
x"20060001",
x"48660003",
x"20030001",
x"08001502",
x"20030000",
x"4860007B",
x"20A70001",
x"A0E30002",
x"4C832800",
x"48BD0003",
x"20030001",
x"E0000000",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08001519",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"0800152F",
x"E8500003",
x"44400006",
x"08001522",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"0800152F",
x"E8300003",
x"44200006",
x"0800152A",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"0800152F",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08001535",
x"20030000",
x"08001537",
x"8CC3FFE8",
x"08001578",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001548",
x"20050001",
x"48650003",
x"20030001",
x"0800154C",
x"20030000",
x"08001578",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"0800156A",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"0800156F",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001574",
x"20050001",
x"48650003",
x"20030001",
x"08001578",
x"20030000",
x"48600003",
x"20E50001",
x"0800148E",
x"20030000",
x"E0000000",
x"20030000",
x"E0000000",
x"A1030002",
x"4C834800",
x"493D0003",
x"20030000",
x"E0000000",
x"A1230002",
x"03E31820",
x"8C660110",
x"C7E1021C",
x"8CC3FFEC",
x"C4600000",
x"44201801",
x"C7E10218",
x"C460FFFC",
x"44202001",
x"C7E10214",
x"C460FFF8",
x"44201001",
x"A1230002",
x"03E31820",
x"8C6703CC",
x"8CC5FFFC",
x"48BC006A",
x"C4E00000",
x"44030001",
x"C4E1FFFC",
x"44010002",
x"C7E502D8",
x"44052802",
x"44A43000",
x"E8D00003",
x"44C02806",
x"080015A1",
x"44C02807",
x"8CC5FFF0",
x"C4A6FFFC",
x"E8A60003",
x"20030000",
x"080015B5",
x"C7E502D4",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"080015AD",
x"44C02807",
x"C4A6FFF8",
x"E8A60003",
x"20030000",
x"080015B5",
x"C8300003",
x"20030001",
x"080015B5",
x"20030000",
x"48600047",
x"C4E0FFF8",
x"44040001",
x"C4E1FFF4",
x"44010002",
x"C7E502DC",
x"44052802",
x"44A33000",
x"E8D00003",
x"44C02806",
x"080015C1",
x"44C02807",
x"C4A60000",
x"E8A60003",
x"20030000",
x"080015D4",
x"C7E502D4",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"080015CC",
x"44C02807",
x"C4A6FFF8",
x"E8A60003",
x"20030000",
x"080015D4",
x"C8300003",
x"20030001",
x"080015D4",
x"20030000",
x"48600025",
x"C4E0FFF0",
x"44020801",
x"C4E0FFEC",
x"44202802",
x"C7E102DC",
x"44A10802",
x"44231000",
x"E8500003",
x"44400806",
x"080015E0",
x"44400807",
x"C4A20000",
x"E8220003",
x"20030000",
x"080015F3",
x"C7E102D8",
x"44A10802",
x"44241000",
x"E8500003",
x"44400806",
x"080015EB",
x"44400807",
x"C4A2FFFC",
x"E8220003",
x"20030000",
x"080015F3",
x"C8100003",
x"20030001",
x"080015F3",
x"20030000",
x"48600003",
x"20030000",
x"080015F8",
x"E7E50208",
x"20030003",
x"080015FB",
x"E7E00208",
x"20030002",
x"080015FE",
x"E7E00208",
x"20030001",
x"08001652",
x"20030002",
x"48A30010",
x"C4E00000",
x"E8100003",
x"20030000",
x"0800160F",
x"C4E0FFFC",
x"44030802",
x"C4E0FFF8",
x"44040002",
x"44200800",
x"C4E0FFF4",
x"44020002",
x"44200000",
x"E7E00208",
x"20030001",
x"08001652",
x"C4E00000",
x"C8100040",
x"C4E1FFFC",
x"44232802",
x"C4E1FFF8",
x"44240802",
x"44A12800",
x"C4E1FFF4",
x"44220802",
x"44A10800",
x"44633002",
x"8CC3FFF0",
x"C4650000",
x"44C53802",
x"44843002",
x"C465FFFC",
x"44C52802",
x"44E53800",
x"44423002",
x"C465FFF8",
x"44C52802",
x"44E53000",
x"8CC3FFF4",
x"48600003",
x"44C02806",
x"08001637",
x"44823802",
x"8CC3FFDC",
x"C4650000",
x"44E52802",
x"44C53000",
x"44432802",
x"C462FFFC",
x"44A21002",
x"44C23000",
x"44641802",
x"C462FFF8",
x"44622802",
x"44C52800",
x"20030003",
x"48A30003",
x"44B11001",
x"0800163C",
x"44A01006",
x"44211802",
x"44020002",
x"44600001",
x"EA000003",
x"20030000",
x"08001650",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"0800164F",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"08001652",
x"20030000",
x"C7E00208",
x"48600003",
x"20030000",
x"0800165C",
x"2003009C",
x"C4610000",
x"E8010003",
x"20030000",
x"0800165C",
x"20030001",
x"4860000A",
x"A1230002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600003",
x"20030000",
x"E0000000",
x"21080001",
x"0800157F",
x"20030098",
x"C4610000",
x"44010000",
x"C7E10134",
x"44201002",
x"C7E1021C",
x"44412800",
x"C7E10130",
x"44201002",
x"C7E10218",
x"44412000",
x"C7E1012C",
x"44200802",
x"C7E00214",
x"44201800",
x"8C850000",
x"AC240000",
x"48BD0003",
x"20030001",
x"080016F0",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"0800168A",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"080016A0",
x"E8500003",
x"44400006",
x"08001693",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"080016A0",
x"E8300003",
x"44200006",
x"0800169B",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"080016A0",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"080016A6",
x"20030000",
x"080016A8",
x"8CC3FFE8",
x"080016E9",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080016B9",
x"20050001",
x"48650003",
x"20030001",
x"080016BD",
x"20030000",
x"080016E9",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"080016DB",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"080016E0",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080016E5",
x"20050001",
x"48650003",
x"20030001",
x"080016E9",
x"20030000",
x"48600006",
x"20050001",
x"40210008",
x"C000148E",
x"20210008",
x"080016F0",
x"20030000",
x"48600004",
x"21080001",
x"8C240000",
x"0800157F",
x"20030001",
x"E0000000",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600073",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600063",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600053",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600043",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600033",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600023",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600013",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C000157F",
x"20210004",
x"48600003",
x"216B0001",
x"080016F6",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"A1830002",
x"4DA35000",
x"8D440000",
x"489D0003",
x"20030000",
x"E0000000",
x"20030063",
x"AC2A0000",
x"48830003",
x"20030001",
x"080018C3",
x"A0830002",
x"03E31820",
x"8C650110",
x"C7E1021C",
x"8CA3FFEC",
x"C4600000",
x"44201801",
x"C7E10218",
x"C460FFFC",
x"44202001",
x"C7E10214",
x"C460FFF8",
x"44200801",
x"A0830002",
x"03E31820",
x"8C6603CC",
x"8CA4FFFC",
x"489C006A",
x"C4C00000",
x"44031001",
x"C4C0FFFC",
x"44403002",
x"C7E202D8",
x"44C21002",
x"44442800",
x"E8B00003",
x"44A01006",
x"0800179F",
x"44A01007",
x"8CA4FFF0",
x"C485FFFC",
x"E8450003",
x"20030000",
x"080017B3",
x"C7E202D4",
x"44C21002",
x"44412800",
x"E8B00003",
x"44A01006",
x"080017AB",
x"44A01007",
x"C485FFF8",
x"E8450003",
x"20030000",
x"080017B3",
x"C8100003",
x"20030001",
x"080017B3",
x"20030000",
x"48600047",
x"C4C0FFF8",
x"44040001",
x"C4C6FFF4",
x"44062802",
x"C7E002DC",
x"44A00002",
x"44031000",
x"E8500003",
x"44400006",
x"080017BF",
x"44400007",
x"C4820000",
x"E8020003",
x"20030000",
x"080017D2",
x"C7E002D4",
x"44A00002",
x"44011000",
x"E8500003",
x"44400006",
x"080017CA",
x"44400007",
x"C482FFF8",
x"E8020003",
x"20030000",
x"080017D2",
x"C8D00003",
x"20030001",
x"080017D2",
x"20030000",
x"48600025",
x"C4C0FFF0",
x"44010001",
x"C4C5FFEC",
x"44051002",
x"C7E002DC",
x"44400002",
x"44030800",
x"E8300003",
x"44200006",
x"080017DE",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"080017F1",
x"C7E002D8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"080017E9",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"080017F1",
x"C8B00003",
x"20030001",
x"080017F1",
x"20030000",
x"48600003",
x"20030000",
x"080017F6",
x"E7E20208",
x"20030003",
x"080017F9",
x"E7E50208",
x"20030002",
x"080017FC",
x"E7E60208",
x"20030001",
x"08001850",
x"20030002",
x"48830010",
x"C4C00000",
x"E8100003",
x"20030000",
x"0800180D",
x"C4C0FFFC",
x"44031002",
x"C4C0FFF8",
x"44040002",
x"44401000",
x"C4C0FFF4",
x"44010002",
x"44400000",
x"E7E00208",
x"20030001",
x"08001850",
x"C4C00000",
x"C8100040",
x"C4C2FFFC",
x"44432802",
x"C4C2FFF8",
x"44441002",
x"44A22800",
x"C4C2FFF4",
x"44411002",
x"44A21000",
x"44633002",
x"8CA3FFF0",
x"C4650000",
x"44C53802",
x"44843002",
x"C465FFFC",
x"44C52802",
x"44E53800",
x"44213002",
x"C465FFF8",
x"44C52802",
x"44E53000",
x"8CA3FFF4",
x"48600003",
x"44C02806",
x"08001835",
x"44813802",
x"8CA3FFDC",
x"C4650000",
x"44E52802",
x"44C53000",
x"44232802",
x"C461FFFC",
x"44A10802",
x"44C13000",
x"44641802",
x"C461FFF8",
x"44612802",
x"44C52800",
x"20030003",
x"48830003",
x"44B10801",
x"0800183A",
x"44A00806",
x"44421802",
x"44010002",
x"44600001",
x"EA000003",
x"20030000",
x"0800184E",
x"8CA3FFE8",
x"48600007",
x"44000004",
x"44400801",
x"C4C0FFF0",
x"44200002",
x"E7E00208",
x"0800184D",
x"44000004",
x"44400800",
x"C4C0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"08001850",
x"20030000",
x"48600003",
x"20030000",
x"080018C3",
x"C7E10208",
x"20030094",
x"C4600000",
x"E8200003",
x"20030000",
x"080018C3",
x"8D44FFFC",
x"489D0003",
x"20030000",
x"080018BF",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860005A",
x"8D44FFF8",
x"489D0003",
x"20030000",
x"080018BD",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860004C",
x"8D44FFF4",
x"489D0003",
x"20030000",
x"080018BB",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860003E",
x"8D44FFF0",
x"489D0003",
x"20030000",
x"080018B9",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600030",
x"8D44FFEC",
x"489D0003",
x"20030000",
x"080018B7",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600022",
x"8D44FFE8",
x"489D0003",
x"20030000",
x"080018B5",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600014",
x"8D44FFE4",
x"489D0003",
x"20030000",
x"080018B3",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600006",
x"200B0008",
x"40210008",
x"C00016F6",
x"20210008",
x"080018B3",
x"20030001",
x"080018B5",
x"20030001",
x"080018B7",
x"20030001",
x"080018B9",
x"20030001",
x"080018BB",
x"20030001",
x"080018BD",
x"20030001",
x"080018BF",
x"20030001",
x"48600003",
x"20030000",
x"080018C3",
x"20030001",
x"48600003",
x"218C0001",
x"08001777",
x"8C2A0000",
x"8D44FFFC",
x"489D0003",
x"20030000",
x"0800192D",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860005A",
x"8D44FFF8",
x"489D0003",
x"20030000",
x"0800192B",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860004C",
x"8D44FFF4",
x"489D0003",
x"20030000",
x"08001929",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"4860003E",
x"8D44FFF0",
x"489D0003",
x"20030000",
x"08001927",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600030",
x"8D44FFEC",
x"489D0003",
x"20030000",
x"08001925",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600022",
x"8D44FFE8",
x"489D0003",
x"20030000",
x"08001923",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600014",
x"8D44FFE4",
x"489D0003",
x"20030000",
x"08001921",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C000157F",
x"20210008",
x"48600006",
x"200B0008",
x"40210008",
x"C00016F6",
x"20210008",
x"08001921",
x"20030001",
x"08001923",
x"20030001",
x"08001925",
x"20030001",
x"08001927",
x"20030001",
x"08001929",
x"20030001",
x"0800192B",
x"20030001",
x"0800192D",
x"20030001",
x"48600003",
x"218C0001",
x"08001777",
x"20030001",
x"E0000000",
x"A1630002",
x"4C835000",
x"495D0002",
x"E0000000",
x"A1430002",
x"03E31820",
x"8C670110",
x"C7E10270",
x"8CE3FFEC",
x"C4600000",
x"44203001",
x"C7E1026C",
x"C460FFFC",
x"44203801",
x"C7E10268",
x"C460FFF8",
x"44202801",
x"8CE3FFFC",
x"487C0087",
x"C5220000",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"0800194D",
x"20060001",
x"C4A10000",
x"48660003",
x"44200007",
x"08001952",
x"44200006",
x"44060001",
x"44021003",
x"C520FFFC",
x"44400002",
x"44070800",
x"E8300003",
x"44200006",
x"0800195B",
x"44200007",
x"C4A1FFFC",
x"E8010003",
x"20080000",
x"0800196C",
x"C520FFF8",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08001966",
x"44200007",
x"C4A1FFF8",
x"E8010003",
x"20080000",
x"0800196C",
x"E7E20208",
x"20080001",
x"0800196E",
x"20080000",
x"4900005B",
x"C522FFFC",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"08001977",
x"20060001",
x"C4A1FFFC",
x"48660003",
x"44200007",
x"0800197C",
x"44200006",
x"44070001",
x"44021003",
x"C520FFF8",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08001985",
x"44200007",
x"C4A1FFF8",
x"E8010003",
x"20080000",
x"08001996",
x"C5200000",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"08001990",
x"44200007",
x"C4A10000",
x"E8010003",
x"20080000",
x"08001996",
x"E7E20208",
x"20080001",
x"08001998",
x"20080000",
x"4900002F",
x"C522FFF8",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"080019A1",
x"20060001",
x"C4A1FFF8",
x"48660003",
x"44200007",
x"080019A6",
x"44200006",
x"44050001",
x"44021003",
x"C5200000",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"080019AF",
x"44200007",
x"C4A10000",
x"E8010003",
x"20080000",
x"080019C0",
x"C520FFFC",
x"44400002",
x"44070800",
x"E8300003",
x"44200006",
x"080019BA",
x"44200007",
x"C4A1FFFC",
x"E8010003",
x"20080000",
x"080019C0",
x"E7E20208",
x"20080001",
x"080019C2",
x"20080000",
x"49000003",
x"20080000",
x"080019C6",
x"20080003",
x"080019C8",
x"20080002",
x"080019CA",
x"20080001",
x"08001A55",
x"20080002",
x"4868001A",
x"8CE3FFF0",
x"C5200000",
x"C4640000",
x"44040802",
x"C520FFFC",
x"C463FFFC",
x"44030002",
x"44201000",
x"C520FFF8",
x"C461FFF8",
x"44010002",
x"44400000",
x"EA000003",
x"20080000",
x"080019E5",
x"44862002",
x"44671002",
x"44821000",
x"44250802",
x"44410800",
x"44200807",
x"44200003",
x"E7E00208",
x"20080001",
x"08001A55",
x"C5210000",
x"C522FFFC",
x"C520FFF8",
x"44211802",
x"8CE5FFF0",
x"C4AA0000",
x"446A2002",
x"44421802",
x"C4ACFFFC",
x"446C1802",
x"44832000",
x"44001802",
x"C4ABFFF8",
x"446B1802",
x"44831800",
x"8CE6FFF4",
x"48C00003",
x"44604806",
x"08001A06",
x"44404002",
x"8CE5FFDC",
x"C4A40000",
x"45042002",
x"44644000",
x"44012002",
x"C4A3FFFC",
x"44831802",
x"45034000",
x"44222002",
x"C4A3FFF8",
x"44834802",
x"45094800",
x"C930004E",
x"44261802",
x"446A2002",
x"44471802",
x"446C1802",
x"44832000",
x"44051802",
x"446B1802",
x"44834000",
x"48C00003",
x"45001806",
x"08001A26",
x"44072002",
x"44451802",
x"44832000",
x"8CE5FFDC",
x"C4A30000",
x"44832002",
x"44251802",
x"44060002",
x"44601800",
x"C4A0FFFC",
x"44600002",
x"44800000",
x"44271802",
x"44460802",
x"44611000",
x"C4A1FFF8",
x"44410802",
x"44010000",
x"44151802",
x"45031800",
x"44C60002",
x"440A0802",
x"44E70002",
x"440C0002",
x"44200800",
x"44A50002",
x"440B0002",
x"44200800",
x"48C00003",
x"44200006",
x"08001A3E",
x"44E51002",
x"8CE5FFDC",
x"C4A00000",
x"44400002",
x"44201000",
x"44A60802",
x"C4A0FFFC",
x"44200002",
x"44401000",
x"44C70802",
x"C4A0FFF8",
x"44200002",
x"44400000",
x"20050003",
x"48650003",
x"44110801",
x"08001A43",
x"44000806",
x"44631002",
x"45210002",
x"44400001",
x"EA000003",
x"20080000",
x"08001A53",
x"44000004",
x"8CE3FFE8",
x"48600003",
x"44000807",
x"08001A4F",
x"44000806",
x"44230001",
x"44090003",
x"E7E00208",
x"20080001",
x"08001A55",
x"20080000",
x"49000009",
x"A1430002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600002",
x"E0000000",
x"216B0001",
x"08001932",
x"C7E00208",
x"AC240000",
x"EA000002",
x"08001AFC",
x"C7E10210",
x"E8010002",
x"08001AFC",
x"20030098",
x"C4610000",
x"44014800",
x"C5200000",
x"44090802",
x"C7E00270",
x"44202800",
x"C520FFFC",
x"44090802",
x"C7E0026C",
x"44202000",
x"C520FFF8",
x"44090802",
x"C7E00268",
x"44201800",
x"8C850000",
x"E4230004",
x"E4240008",
x"E425000C",
x"48BD0003",
x"20030001",
x"08001AF1",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08001A8B",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"08001AA1",
x"E8500003",
x"44400006",
x"08001A94",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"08001AA1",
x"E8300003",
x"44200006",
x"08001A9C",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"08001AA1",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08001AA7",
x"20030000",
x"08001AA9",
x"8CC3FFE8",
x"08001AEA",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001ABA",
x"20050001",
x"48650003",
x"20030001",
x"08001ABE",
x"20030000",
x"08001AEA",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"08001ADC",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"08001AE1",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001AE6",
x"20050001",
x"48650003",
x"20030001",
x"08001AEA",
x"20030000",
x"48600006",
x"20050001",
x"40210014",
x"C000148E",
x"20210014",
x"08001AF1",
x"20030000",
x"48600002",
x"08001AFC",
x"E7E90210",
x"C425000C",
x"E7E5021C",
x"C4240008",
x"E7E40218",
x"C4230004",
x"E7E30214",
x"AFEA0220",
x"AFE8020C",
x"216B0001",
x"8C240000",
x"08001932",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"AC290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"21AD0001",
x"8C290000",
x"08001AFF",
x"A1C30002",
x"4DE36000",
x"8D830000",
x"487D0002",
x"E0000000",
x"20040063",
x"AC290000",
x"48640053",
x"8D83FFFC",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF8",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF4",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF0",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFEC",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFE8",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFE4",
x"487D0002",
x"08001BC2",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"200D0008",
x"8C290000",
x"40210008",
x"C0001AFF",
x"20210008",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C660110",
x"C7E10270",
x"8CC3FFEC",
x"C4600000",
x"44202801",
x"C7E1026C",
x"C460FFFC",
x"44203001",
x"C7E10268",
x"C460FFF8",
x"44202001",
x"8CC4FFFC",
x"489C0087",
x"C5220000",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"08001BDA",
x"20050001",
x"C4810000",
x"48650003",
x"44200007",
x"08001BDF",
x"44200006",
x"44050001",
x"44021003",
x"C520FFFC",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"08001BE8",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"08001BF9",
x"C520FFF8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"08001BF3",
x"44200007",
x"C481FFF8",
x"E8010003",
x"20030000",
x"08001BF9",
x"E7E20208",
x"20030001",
x"08001BFB",
x"20030000",
x"4860005B",
x"C522FFFC",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"08001C04",
x"20050001",
x"C481FFFC",
x"48650003",
x"44200007",
x"08001C09",
x"44200006",
x"44060001",
x"44021003",
x"C520FFF8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"08001C12",
x"44200007",
x"C481FFF8",
x"E8010003",
x"20030000",
x"08001C23",
x"C5200000",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08001C1D",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"08001C23",
x"E7E20208",
x"20030001",
x"08001C25",
x"20030000",
x"4860002F",
x"C522FFF8",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"08001C2E",
x"20050001",
x"C481FFF8",
x"48650003",
x"44200007",
x"08001C33",
x"44200006",
x"44040001",
x"44021003",
x"C5200000",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08001C3C",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"08001C4D",
x"C520FFFC",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"08001C47",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"08001C4D",
x"E7E20208",
x"20030001",
x"08001C4F",
x"20030000",
x"48600003",
x"20030000",
x"08001C53",
x"20030003",
x"08001C55",
x"20030002",
x"08001C57",
x"20030001",
x"08001CE2",
x"20030002",
x"4883001A",
x"8CC3FFF0",
x"C5200000",
x"C4670000",
x"44070802",
x"C520FFFC",
x"C463FFFC",
x"44030002",
x"44201000",
x"C520FFF8",
x"C461FFF8",
x"44010002",
x"44400000",
x"EA000003",
x"20030000",
x"08001C72",
x"44E52802",
x"44661002",
x"44A21000",
x"44240802",
x"44410800",
x"44200807",
x"44200003",
x"E7E00208",
x"20030001",
x"08001CE2",
x"C5210000",
x"C522FFFC",
x"C520FFF8",
x"44211802",
x"8CC3FFF0",
x"C4690000",
x"44693802",
x"44421802",
x"C46BFFFC",
x"446B1802",
x"44E33800",
x"44001802",
x"C46AFFF8",
x"446A1802",
x"44E31800",
x"8CC5FFF4",
x"48A00003",
x"44604006",
x"08001C93",
x"44404002",
x"8CC3FFDC",
x"C4670000",
x"45073802",
x"44674000",
x"44013802",
x"C463FFFC",
x"44E31802",
x"45036000",
x"44223802",
x"C463FFF8",
x"44E34002",
x"45884000",
x"C910004E",
x"44251802",
x"44693802",
x"44461802",
x"446B1802",
x"44E33800",
x"44041802",
x"446A1802",
x"44E33800",
x"48A00003",
x"44E01806",
x"08001CB3",
x"44066002",
x"44441802",
x"45836000",
x"8CC3FFDC",
x"C4630000",
x"45831802",
x"44246002",
x"44050002",
x"45806000",
x"C460FFFC",
x"45800002",
x"44600000",
x"44261802",
x"44450802",
x"44611000",
x"C461FFF8",
x"44410802",
x"44010000",
x"44151802",
x"44E31800",
x"44A50002",
x"44090802",
x"44C60002",
x"440B0002",
x"44200800",
x"44840002",
x"440A0002",
x"44200800",
x"48A00003",
x"44200006",
x"08001CCB",
x"44C41002",
x"8CC3FFDC",
x"C4600000",
x"44400002",
x"44201000",
x"44850802",
x"C460FFFC",
x"44200002",
x"44401000",
x"44A60802",
x"C460FFF8",
x"44200002",
x"44400000",
x"20030003",
x"48830003",
x"44110801",
x"08001CD0",
x"44000806",
x"44631002",
x"45010002",
x"44400001",
x"EA000003",
x"20030000",
x"08001CE0",
x"44000004",
x"8CC3FFE8",
x"48600003",
x"44000807",
x"08001CDC",
x"44000806",
x"44230001",
x"44080003",
x"E7E00208",
x"20030001",
x"08001CE2",
x"20030000",
x"48600002",
x"08001D39",
x"C7E00208",
x"C7E10210",
x"E8010002",
x"08001D39",
x"8D83FFFC",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF8",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF4",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFF0",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFEC",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFE8",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"8D83FFE4",
x"487D0002",
x"08001D39",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C0001932",
x"20210008",
x"200D0008",
x"8C290000",
x"40210008",
x"C0001AFF",
x"20210008",
x"21CE0001",
x"8C290000",
x"08001B69",
x"A1430002",
x"4C834800",
x"493D0002",
x"E0000000",
x"A1230002",
x"03E31820",
x"8C660110",
x"8CC5FFD8",
x"C4A30000",
x"C4A4FFFC",
x"C4A2FFF8",
x"A1230002",
x"4D633800",
x"8CC3FFFC",
x"487C006A",
x"C4E00000",
x"44030001",
x"C4E1FFFC",
x"44010002",
x"C585FFFC",
x"44052802",
x"44A43000",
x"E8D00003",
x"44C02806",
x"08001D56",
x"44C02807",
x"8CC3FFF0",
x"C466FFFC",
x"E8A60003",
x"20080000",
x"08001D6A",
x"C585FFF8",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"08001D62",
x"44C02807",
x"C466FFF8",
x"E8A60003",
x"20080000",
x"08001D6A",
x"C8300003",
x"20080001",
x"08001D6A",
x"20080000",
x"49000047",
x"C4E0FFF8",
x"44040001",
x"C4E1FFF4",
x"44010002",
x"C5850000",
x"44052802",
x"44A33000",
x"E8D00003",
x"44C02806",
x"08001D76",
x"44C02807",
x"C4660000",
x"E8A60003",
x"20080000",
x"08001D89",
x"C585FFF8",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"08001D81",
x"44C02807",
x"C466FFF8",
x"E8A60003",
x"20080000",
x"08001D89",
x"C8300003",
x"20080001",
x"08001D89",
x"20080000",
x"49000025",
x"C4E0FFF0",
x"44020801",
x"C4E0FFEC",
x"44202802",
x"C5810000",
x"44A10802",
x"44231000",
x"E8500003",
x"44400806",
x"08001D95",
x"44400807",
x"C4620000",
x"E8220003",
x"20080000",
x"08001DA8",
x"C581FFFC",
x"44A10802",
x"44241000",
x"E8500003",
x"44400806",
x"08001DA0",
x"44400807",
x"C462FFFC",
x"E8220003",
x"20080000",
x"08001DA8",
x"C8100003",
x"20080001",
x"08001DA8",
x"20080000",
x"49000003",
x"20080000",
x"08001DAD",
x"E7E50208",
x"20080003",
x"08001DB0",
x"E7E00208",
x"20080002",
x"08001DB3",
x"E7E00208",
x"20080001",
x"08001DE0",
x"20080002",
x"4868000A",
x"C4E10000",
x"E8300003",
x"20080000",
x"08001DBE",
x"C4A0FFF4",
x"44200002",
x"E7E00208",
x"20080001",
x"08001DE0",
x"C4E50000",
x"C8B0001F",
x"C4E0FFFC",
x"44030802",
x"C4E0FFF8",
x"44040002",
x"44200800",
x"C4E0FFF4",
x"44020002",
x"44200800",
x"C4A0FFF4",
x"44211002",
x"44A00002",
x"44400001",
x"EA000003",
x"20080000",
x"08001DDE",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"08001DDD",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20080001",
x"08001DE0",
x"20080000",
x"49000009",
x"A1230002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600002",
x"E0000000",
x"214A0001",
x"08001D3C",
x"C7E00208",
x"AC240000",
x"EA000002",
x"08001E87",
x"C7E10210",
x"E8010002",
x"08001E87",
x"20030098",
x"C4610000",
x"44014800",
x"C5800000",
x"44090802",
x"C7E0027C",
x"44202800",
x"C580FFFC",
x"44090802",
x"C7E00278",
x"44202000",
x"C580FFF8",
x"44090802",
x"C7E00274",
x"44201800",
x"8C850000",
x"E4230004",
x"E4240008",
x"E425000C",
x"48BD0003",
x"20030001",
x"08001E7C",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08001E16",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"08001E2C",
x"E8500003",
x"44400006",
x"08001E1F",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"08001E2C",
x"E8300003",
x"44200006",
x"08001E27",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"08001E2C",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08001E32",
x"20030000",
x"08001E34",
x"8CC3FFE8",
x"08001E75",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001E45",
x"20050001",
x"48650003",
x"20030001",
x"08001E49",
x"20030000",
x"08001E75",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"08001E67",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"08001E6C",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001E71",
x"20050001",
x"48650003",
x"20030001",
x"08001E75",
x"20030000",
x"48600006",
x"20050001",
x"40210014",
x"C000148E",
x"20210014",
x"08001E7C",
x"20030000",
x"48600002",
x"08001E87",
x"E7E90210",
x"C425000C",
x"E7E5021C",
x"C4240008",
x"E7E40218",
x"C4230004",
x"E7E30214",
x"AFE90220",
x"AFE8020C",
x"214A0001",
x"8C240000",
x"08001D3C",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"22100001",
x"08001E8A",
x"A2630002",
x"4E837800",
x"8DE30000",
x"487D0002",
x"E0000000",
x"20040063",
x"4864005A",
x"8DE3FFFC",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF8",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF4",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF0",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFEC",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFE8",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFE4",
x"487D0002",
x"08001F5A",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20100008",
x"222D0000",
x"224E0000",
x"C0001E8A",
x"20210004",
x"08002059",
x"A0640002",
x"03E42020",
x"8C860110",
x"8CC5FFD8",
x"C4A20000",
x"C4A3FFFC",
x"C4A1FFF8",
x"A0630002",
x"4E233800",
x"8CC4FFFC",
x"489C006A",
x"C4E00000",
x"44022001",
x"C4E0FFFC",
x"44803002",
x"C644FFFC",
x"44C42002",
x"44832800",
x"E8B00003",
x"44A02006",
x"08001F71",
x"44A02007",
x"8CC4FFF0",
x"C485FFFC",
x"E8850003",
x"20030000",
x"08001F85",
x"C644FFF8",
x"44C42002",
x"44812800",
x"E8B00003",
x"44A02006",
x"08001F7D",
x"44A02007",
x"C485FFF8",
x"E8850003",
x"20030000",
x"08001F85",
x"C8100003",
x"20030001",
x"08001F85",
x"20030000",
x"48600047",
x"C4E0FFF8",
x"44030001",
x"C4E6FFF4",
x"44062802",
x"C6400000",
x"44A00002",
x"44022000",
x"E8900003",
x"44800006",
x"08001F91",
x"44800007",
x"C4840000",
x"E8040003",
x"20030000",
x"08001FA4",
x"C640FFF8",
x"44A00002",
x"44012000",
x"E8900003",
x"44800006",
x"08001F9C",
x"44800007",
x"C484FFF8",
x"E8040003",
x"20030000",
x"08001FA4",
x"C8D00003",
x"20030001",
x"08001FA4",
x"20030000",
x"48600025",
x"C4E0FFF0",
x"44010001",
x"C4E5FFEC",
x"44052002",
x"C6400000",
x"44800002",
x"44020800",
x"E8300003",
x"44200006",
x"08001FB0",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"08001FC3",
x"C640FFFC",
x"44800002",
x"44030800",
x"E8300003",
x"44200006",
x"08001FBB",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"08001FC3",
x"C8B00003",
x"20030001",
x"08001FC3",
x"20030000",
x"48600003",
x"20030000",
x"08001FC8",
x"E7E40208",
x"20030003",
x"08001FCB",
x"E7E50208",
x"20030002",
x"08001FCE",
x"E7E60208",
x"20030001",
x"08001FFB",
x"20030002",
x"4883000A",
x"C4E10000",
x"E8300003",
x"20030000",
x"08001FD9",
x"C4A0FFF4",
x"44200002",
x"E7E00208",
x"20030001",
x"08001FFB",
x"C4E40000",
x"C890001F",
x"C4E0FFFC",
x"44021002",
x"C4E0FFF8",
x"44030002",
x"44401000",
x"C4E0FFF4",
x"44010002",
x"44400800",
x"C4A0FFF4",
x"44211002",
x"44800002",
x"44400001",
x"EA000003",
x"20030000",
x"08001FF9",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"08001FF8",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"08001FFB",
x"20030000",
x"48600002",
x"08002059",
x"C7E00208",
x"C7E10210",
x"E8010002",
x"08002059",
x"8DE3FFFC",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF8",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF4",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFF0",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFEC",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFE8",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20210004",
x"8DE3FFE4",
x"487D0002",
x"08002059",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0001D3C",
x"20100008",
x"222D0000",
x"224E0000",
x"C0001E8A",
x"20210004",
x"22730001",
x"08001EFB",
x"6AA00064",
x"A2A30002",
x"03E31820",
x"8C7706B4",
x"8EF8FFFC",
x"200300D4",
x"C4600000",
x"E7E00210",
x"20130000",
x"8FF40204",
x"8F11FFFC",
x"8F120000",
x"40210004",
x"C0001EFB",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"08002076",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"08002076",
x"20030001",
x"48600002",
x"080020BD",
x"8FE30220",
x"A0640002",
x"8FE3020C",
x"00831820",
x"8EE40000",
x"48640040",
x"200C0000",
x"8FED0204",
x"40210004",
x"C0001777",
x"20210004",
x"48600039",
x"8F030000",
x"C7E0022C",
x"C4620000",
x"44020802",
x"C7E00228",
x"C464FFFC",
x"44040002",
x"44200800",
x"C7E00224",
x"C463FFF8",
x"44030002",
x"44200800",
x"C6E0FFF8",
x"440B2802",
x"44A10802",
x"C6C50000",
x"44A22802",
x"C6C2FFFC",
x"44441002",
x"44A22000",
x"C6C2FFF8",
x"44431002",
x"44821000",
x"44020002",
x"EA010002",
x"080020AD",
x"C7E30250",
x"C7E20238",
x"44221002",
x"44621000",
x"E7E20250",
x"C7E3024C",
x"C7E20234",
x"44221002",
x"44621000",
x"E7E2024C",
x"C7E30248",
x"C7E20230",
x"44220802",
x"44610800",
x"E7E10248",
x"EA000002",
x"080020BB",
x"44000002",
x"44000002",
x"440A0002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"080020BC",
x"080020BD",
x"42B50001",
x"0800205B",
x"E0000000",
x"20030004",
x"68790415",
x"200300D4",
x"C4600000",
x"E7E00210",
x"200E0000",
x"8FEF0204",
x"22C90000",
x"40210004",
x"C0001B69",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"080020D7",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"080020D7",
x"20030001",
x"48600023",
x"2004FFFF",
x"A3230002",
x"6E632000",
x"4B200002",
x"E0000000",
x"C6C10000",
x"C7E00134",
x"44201002",
x"C6C1FFFC",
x"C7E00130",
x"44200002",
x"44401000",
x"C6C1FFF8",
x"C7E0012C",
x"44200002",
x"44400000",
x"44000007",
x"EA000002",
x"E0000000",
x"44000802",
x"44200002",
x"440D0802",
x"C7E00138",
x"44200002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"E0000000",
x"8FE70220",
x"A0E30002",
x"03E31820",
x"8C630110",
x"8C7EFFF8",
x"8C7AFFE4",
x"C7400000",
x"440D5802",
x"8C64FFFC",
x"489C0016",
x"8FE4020C",
x"E7F0022C",
x"E7F00228",
x"E7F00224",
x"40850001",
x"A0A40002",
x"02C40831",
x"C8300008",
x"EA010004",
x"200400A0",
x"C4800000",
x"08002112",
x"200400C8",
x"C4800000",
x"08002114",
x"46000006",
x"44000007",
x"A0A40002",
x"03E42020",
x"E480022C",
x"08002170",
x"20050002",
x"4885000C",
x"8C64FFF0",
x"C4800000",
x"44000007",
x"E7E0022C",
x"C480FFFC",
x"44000007",
x"E7E00228",
x"C480FFF8",
x"44000007",
x"E7E00224",
x"08002170",
x"C7E1021C",
x"8C64FFEC",
x"C4800000",
x"44202001",
x"C7E10218",
x"C480FFFC",
x"44201801",
x"C7E10214",
x"C480FFF8",
x"44200001",
x"8C64FFF0",
x"C4810000",
x"44810802",
x"C482FFFC",
x"44622802",
x"C482FFF8",
x"44023802",
x"8C64FFF4",
x"48800005",
x"E7E1022C",
x"E7E50228",
x"E7E70224",
x"08002156",
x"8C64FFDC",
x"C482FFF8",
x"44623002",
x"C482FFFC",
x"44021002",
x"44C21000",
x"44551002",
x"44220800",
x"E7E1022C",
x"C481FFF8",
x"44811002",
x"C4810000",
x"44010002",
x"44400000",
x"44150002",
x"44A00000",
x"E7E00228",
x"C480FFFC",
x"44800802",
x"C4800000",
x"44600002",
x"44200000",
x"44150002",
x"44E00000",
x"E7E00224",
x"8C64FFE8",
x"C7E2022C",
x"44420802",
x"C7E00228",
x"44000002",
x"44200800",
x"C7E00224",
x"44000002",
x"44200000",
x"44000804",
x"C8300006",
x"48800003",
x"46210003",
x"08002165",
x"46810003",
x"08002168",
x"200400C8",
x"C4800000",
x"44400802",
x"E7E1022C",
x"C7E10228",
x"44200802",
x"E7E10228",
x"C7E10224",
x"44200002",
x"E7E00224",
x"C7E0021C",
x"E7E00270",
x"C7E00218",
x"E7E0026C",
x"C7E00214",
x"E7E00268",
x"8C640000",
x"8C65FFE0",
x"C4A00000",
x"E7E00238",
x"C4A0FFFC",
x"E7E00234",
x"C4A0FFF8",
x"E7E00230",
x"489C0028",
x"C7E1021C",
x"8C65FFEC",
x"C4A00000",
x"44202801",
x"2003002C",
x"C4690000",
x"44A90002",
x"40210004",
x"C0000051",
x"20030028",
x"C4660000",
x"44060002",
x"44A04001",
x"20030034",
x"C4650000",
x"C7E10214",
x"C4A0FFF8",
x"44203801",
x"44E90002",
x"C0000051",
x"20210004",
x"44060002",
x"44E00801",
x"E9050008",
x"E8250004",
x"200300D8",
x"C4600000",
x"0800219D",
x"200300DC",
x"C4600000",
x"080021A4",
x"E8250004",
x"200300DC",
x"C4600000",
x"080021A4",
x"200300D8",
x"C4600000",
x"E7E00234",
x"080023C0",
x"20050002",
x"48850082",
x"C7E10218",
x"20030030",
x"C4600000",
x"44201002",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"080021B4",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080021DA",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080021CB",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080021C6",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080021CB",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080021DA",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080021D5",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080021DA",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080021FD",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080021EE",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080021E9",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080021EE",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080021FD",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080021F8",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080021FD",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"E8600006",
x"EA020003",
x"20030000",
x"08002202",
x"20030001",
x"08002207",
x"EA020003",
x"20030001",
x"08002207",
x"20030000",
x"E8600003",
x"44000806",
x"0800220B",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800220F",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"08002222",
x"44000806",
x"44210002",
x"47600802",
x"E7E10238",
x"46200001",
x"47600002",
x"E7E00234",
x"080023C0",
x"20050003",
x"48850095",
x"C7E1021C",
x"8C63FFEC",
x"C4600000",
x"44200001",
x"C7E20214",
x"C461FFF8",
x"44410801",
x"44000002",
x"44210802",
x"44010000",
x"44000004",
x"20030034",
x"C4610000",
x"44010003",
x"E4200000",
x"40210008",
x"C0000051",
x"20210008",
x"44000806",
x"C4200000",
x"44010001",
x"441E0002",
x"46C01001",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"0800224A",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08002270",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002261",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800225C",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"08002261",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"08002270",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800226B",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"08002270",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"08002293",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002284",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800227F",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"08002284",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"08002293",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800228E",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"08002293",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"E8600006",
x"EA020003",
x"20030000",
x"08002298",
x"20030001",
x"0800229D",
x"EA020003",
x"20030001",
x"0800229D",
x"20030000",
x"E8600003",
x"44000806",
x"080022A1",
x"47A00801",
x"EAC10003",
x"44200006",
x"080022A5",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"080022B8",
x"44000806",
x"44210002",
x"441B0802",
x"E7E10234",
x"46200001",
x"441B0002",
x"E7E00230",
x"080023C0",
x"20050004",
x"48850100",
x"C7E1021C",
x"8C66FFEC",
x"C4C00000",
x"44200801",
x"8C65FFF0",
x"C4A00000",
x"44000004",
x"44200802",
x"C7E20214",
x"C4C0FFF8",
x"44401001",
x"C4A0FFF8",
x"44000004",
x"44401002",
x"44211802",
x"44420002",
x"44602800",
x"E8300003",
x"44200006",
x"080022D6",
x"44200007",
x"2003008C",
x"C4660000",
x"E806005D",
x"44410803",
x"E8300003",
x"44200006",
x"080022DE",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"080022E3",
x"2003FFFF",
x"080022E5",
x"20030001",
x"48600003",
x"44001806",
x"080022E9",
x"46201803",
x"44630002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44202002",
x"20040078",
x"C4810000",
x"44220800",
x"44811003",
x"20040074",
x"C4810000",
x"44202002",
x"20040070",
x"C4810000",
x"44220800",
x"44811003",
x"2004006C",
x"C4810000",
x"44202002",
x"20040068",
x"C4810000",
x"44220800",
x"44811003",
x"20040064",
x"C4810000",
x"44202002",
x"47820800",
x"44811003",
x"20040060",
x"C4810000",
x"44202002",
x"2004005C",
x"C4810000",
x"44220800",
x"44811003",
x"20040058",
x"C4810000",
x"44202002",
x"20040054",
x"C4810000",
x"44220800",
x"44811003",
x"20040050",
x"C4810000",
x"44202002",
x"47220800",
x"44810803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44202002",
x"47020800",
x"44810803",
x"46E10800",
x"44010003",
x"46200000",
x"44600803",
x"68030006",
x"68600003",
x"44200006",
x"0800232E",
x"47E10001",
x"08002330",
x"46C10001",
x"20030044",
x"C4610000",
x"44010002",
x"441E0003",
x"08002337",
x"20030088",
x"C4600000",
x"E4200004",
x"4021000C",
x"C0000051",
x"2021000C",
x"44000806",
x"C4200004",
x"44013801",
x"C7E10218",
x"C4C0FFFC",
x"44200801",
x"C4A0FFFC",
x"44000004",
x"44200802",
x"E8B00003",
x"44A00006",
x"08002348",
x"44A00007",
x"E806005D",
x"44250803",
x"E8300003",
x"44200006",
x"0800234E",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"08002353",
x"2003FFFF",
x"08002355",
x"20030001",
x"48600003",
x"44002006",
x"08002359",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44610803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800003",
x"68030006",
x"68600003",
x"44000806",
x"0800239E",
x"47E00801",
x"080023A0",
x"46C00801",
x"20030044",
x"C4600000",
x"44200002",
x"441E0003",
x"080023A7",
x"20030088",
x"C4600000",
x"E4200008",
x"40210010",
x"C0000051",
x"20210010",
x"44000806",
x"C4200008",
x"44010001",
x"2003003C",
x"C4620000",
x"46A70801",
x"44210802",
x"44410801",
x"46A00001",
x"44000002",
x"44200801",
x"E8300003",
x"44200006",
x"080023BA",
x"46000006",
x"47600802",
x"20030038",
x"C4600000",
x"44200003",
x"E7E00230",
x"080023C0",
x"A0E40002",
x"8FE3020C",
x"00832020",
x"A3230002",
x"6E632000",
x"A3230002",
x"4E831800",
x"C7E0021C",
x"E4600000",
x"C7E00218",
x"E460FFFC",
x"C7E00214",
x"E460FFF8",
x"C7400000",
x"E8150023",
x"20040001",
x"A3230002",
x"6E432000",
x"A3230002",
x"4E231800",
x"C7E00238",
x"E4600000",
x"C7E00234",
x"E460FFFC",
x"C7E00230",
x"E460FFF8",
x"A3230002",
x"4E232000",
x"20030024",
x"C4600000",
x"440B0002",
x"C4810000",
x"44200802",
x"E4810000",
x"C481FFFC",
x"44200802",
x"E481FFFC",
x"C481FFF8",
x"44200002",
x"E480FFF8",
x"A3230002",
x"4E031800",
x"C7E0022C",
x"E4600000",
x"C7E00228",
x"E460FFFC",
x"C7E00224",
x"E460FFF8",
x"080023F4",
x"20040000",
x"A3230002",
x"6E432000",
x"20030020",
x"C4630000",
x"C6C10000",
x"C7E0022C",
x"44202802",
x"C6C4FFFC",
x"C7E20228",
x"44821002",
x"44A22800",
x"C6C4FFF8",
x"C7E20224",
x"44821002",
x"44A21000",
x"44621002",
x"44400002",
x"44200000",
x"E6C00000",
x"C6C1FFFC",
x"C7E00228",
x"44400002",
x"44200000",
x"E6C0FFFC",
x"C6C1FFF8",
x"C7E00224",
x"44400002",
x"44200000",
x"E6C0FFF8",
x"C740FFFC",
x"45A05002",
x"200C0000",
x"8FED0204",
x"40210010",
x"C0001777",
x"20210010",
x"48600037",
x"C7E1022C",
x"C7E00134",
x"44201002",
x"C7E10228",
x"C7E30130",
x"44230802",
x"44412000",
x"C7E10224",
x"C7E2012C",
x"44220802",
x"44810800",
x"44200807",
x"442B0802",
x"C6C40000",
x"44802002",
x"C6C0FFFC",
x"44030002",
x"44801800",
x"C6C0FFF8",
x"44020002",
x"44600000",
x"44000007",
x"EA010002",
x"0800243E",
x"C7E30250",
x"C7E20238",
x"44221002",
x"44621000",
x"E7E20250",
x"C7E3024C",
x"C7E20234",
x"44221002",
x"44621000",
x"E7E2024C",
x"C7E30248",
x"C7E20230",
x"44220802",
x"44610800",
x"E7E10248",
x"EA000002",
x"0800244C",
x"44000002",
x"44000002",
x"440A0002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"0800244D",
x"C7E0021C",
x"E7E0027C",
x"C7E00218",
x"E7E00278",
x"C7E00214",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7E1021C",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C7E10218",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C7E10214",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"080024A1",
x"20050002",
x"68A60002",
x"080024A1",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"0800249B",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"080024A0",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"43E3021C",
x"40210010",
x"C00013F1",
x"20210010",
x"080024A7",
x"8FE306B8",
x"40630001",
x"AC36000C",
x"AC300010",
x"AC350014",
x"AC370018",
x"AC31001C",
x"AC320020",
x"AC330024",
x"AC340028",
x"AC38002C",
x"AC330030",
x"20750000",
x"40210038",
x"C000205B",
x"20210038",
x"200300A4",
x"C4600000",
x"E80D0002",
x"E0000000",
x"20030004",
x"6B230002",
x"080024C3",
x"23230001",
x"2004FFFF",
x"A0630002",
x"8C330030",
x"6E632000",
x"20030002",
x"4BC30011",
x"C7400000",
x"46200001",
x"45A06802",
x"23390001",
x"C7E00210",
x"45C07000",
x"8C38002C",
x"8C340028",
x"8C330024",
x"8C320020",
x"8C31001C",
x"8C370018",
x"8C350014",
x"8C300010",
x"8C36000C",
x"080020C0",
x"E0000000",
x"E0000000",
x"200400D4",
x"C4800000",
x"E7E00210",
x"20130000",
x"8FF40204",
x"20710000",
x"22B20000",
x"40210004",
x"C0001EFB",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"080024ED",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"080024ED",
x"20030001",
x"48600002",
x"E0000000",
x"8FE30220",
x"A0630002",
x"03E31820",
x"8C6E0110",
x"8DC3FFFC",
x"487C0016",
x"8FE3020C",
x"E7F0022C",
x"E7F00228",
x"E7F00224",
x"40640001",
x"A0830002",
x"02A30831",
x"C8300008",
x"EA010004",
x"200300A0",
x"C4600000",
x"08002503",
x"200300C8",
x"C4600000",
x"08002505",
x"46000006",
x"44000007",
x"A0830002",
x"03E31820",
x"E460022C",
x"08002561",
x"20040002",
x"4864000C",
x"8DC3FFF0",
x"C4600000",
x"44000007",
x"E7E0022C",
x"C460FFFC",
x"44000007",
x"E7E00228",
x"C460FFF8",
x"44000007",
x"E7E00224",
x"08002561",
x"C7E1021C",
x"8DC3FFEC",
x"C4600000",
x"44202001",
x"C7E10218",
x"C460FFFC",
x"44201801",
x"C7E10214",
x"C460FFF8",
x"44200001",
x"8DC3FFF0",
x"C4610000",
x"44811002",
x"C461FFFC",
x"44613002",
x"C461FFF8",
x"44013802",
x"8DC3FFF4",
x"48600005",
x"E7E2022C",
x"E7E60228",
x"E7E70224",
x"08002547",
x"8DC3FFDC",
x"C461FFF8",
x"44612802",
x"C461FFFC",
x"44010802",
x"44A10800",
x"44350802",
x"44410800",
x"E7E1022C",
x"C461FFF8",
x"44811002",
x"C4610000",
x"44010002",
x"44400000",
x"44150002",
x"44C00000",
x"E7E00228",
x"C460FFFC",
x"44800802",
x"C4600000",
x"44600002",
x"44200000",
x"44150002",
x"44E00000",
x"E7E00224",
x"8DC3FFE8",
x"C7E2022C",
x"44420802",
x"C7E00228",
x"44000002",
x"44200800",
x"C7E00224",
x"44000002",
x"44200000",
x"44000804",
x"C8300006",
x"48600003",
x"46210003",
x"08002556",
x"46810003",
x"08002559",
x"200300C8",
x"C4600000",
x"44400802",
x"E7E1022C",
x"C7E10228",
x"44200802",
x"E7E10228",
x"C7E10224",
x"44200002",
x"E7E00224",
x"8DC30000",
x"8DC4FFE0",
x"C4800000",
x"E7E00238",
x"C480FFFC",
x"E7E00234",
x"C480FFF8",
x"E7E00230",
x"487C0028",
x"C7E1021C",
x"8DC5FFEC",
x"C4A00000",
x"44202801",
x"2003002C",
x"C4690000",
x"44A90002",
x"40210004",
x"C0000051",
x"20030028",
x"C4680000",
x"44080002",
x"44A03801",
x"20030034",
x"C4660000",
x"C7E10214",
x"C4A0FFF8",
x"44202801",
x"44A90002",
x"C0000051",
x"20210004",
x"44080002",
x"44A00801",
x"E8E60008",
x"E8260004",
x"200300D8",
x"C4600000",
x"08002588",
x"200300DC",
x"C4600000",
x"0800258F",
x"E8260004",
x"200300DC",
x"C4600000",
x"0800258F",
x"200300D8",
x"C4600000",
x"E7E00234",
x"080027AB",
x"20040002",
x"48640082",
x"C7E10218",
x"20030030",
x"C4600000",
x"44201002",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"0800259F",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080025C5",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080025B6",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080025B1",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080025B6",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080025C5",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080025C0",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080025C5",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080025E8",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080025D9",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080025D4",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080025D9",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"080025E8",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080025E3",
x"443D0800",
x"40210004",
x"C0000A77",
x"20210004",
x"080025E8",
x"443D0801",
x"40210004",
x"C0000A77",
x"20210004",
x"E8600006",
x"EA020003",
x"20030000",
x"080025ED",
x"20030001",
x"080025F2",
x"EA020003",
x"20030001",
x"080025F2",
x"20030000",
x"E8600003",
x"44000806",
x"080025F6",
x"47A00801",
x"EAC10003",
x"44200006",
x"080025FA",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"0800260D",
x"44000806",
x"44210002",
x"47600802",
x"E7E10238",
x"46200001",
x"47600002",
x"E7E00234",
x"080027AB",
x"20040003",
x"48640095",
x"C7E1021C",
x"8DC3FFEC",
x"C4600000",
x"44200801",
x"C7E20214",
x"C460FFF8",
x"44400001",
x"44210802",
x"44000002",
x"44200000",
x"44000004",
x"20030034",
x"C4610000",
x"44010003",
x"E4200000",
x"40210008",
x"C0000051",
x"20210008",
x"44000806",
x"C4200000",
x"44010001",
x"441E0002",
x"46C01001",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"08002635",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"0800265B",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800264C",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002647",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"0800264C",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"0800265B",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002656",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"0800265B",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"0800267E",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800266F",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800266A",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"0800266F",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"0800267E",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002679",
x"443D0800",
x"40210008",
x"C0000A77",
x"20210008",
x"0800267E",
x"443D0801",
x"40210008",
x"C0000A77",
x"20210008",
x"E8600006",
x"EA020003",
x"20030000",
x"08002683",
x"20030001",
x"08002688",
x"EA020003",
x"20030001",
x"08002688",
x"20030000",
x"E8600003",
x"44000806",
x"0800268C",
x"47A00801",
x"EAC10003",
x"44200006",
x"08002690",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"080026A3",
x"44000806",
x"44210002",
x"441B0802",
x"E7E10234",
x"46200001",
x"441B0002",
x"E7E00230",
x"080027AB",
x"20040004",
x"48640100",
x"C7E1021C",
x"8DC5FFEC",
x"C4A00000",
x"44200801",
x"8DC6FFF0",
x"C4C00000",
x"44000004",
x"44200802",
x"C7E20214",
x"C4A0FFF8",
x"44401001",
x"C4C0FFF8",
x"44000004",
x"44401002",
x"44211802",
x"44420002",
x"44602800",
x"E8300003",
x"44200006",
x"080026C1",
x"44200007",
x"2003008C",
x"C4660000",
x"E806005D",
x"44410803",
x"E8300003",
x"44200006",
x"080026C9",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"080026CE",
x"2003FFFF",
x"080026D0",
x"20030001",
x"48600003",
x"44002006",
x"080026D4",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44610803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800803",
x"68030006",
x"68600003",
x"44200006",
x"08002719",
x"47E10001",
x"0800271B",
x"46C10001",
x"20030044",
x"C4610000",
x"44010002",
x"441E0003",
x"08002722",
x"20030088",
x"C4600000",
x"E4200004",
x"4021000C",
x"C0000051",
x"2021000C",
x"44000806",
x"C4200004",
x"44013801",
x"C7E10218",
x"C4A0FFFC",
x"44200801",
x"C4C0FFFC",
x"44000004",
x"44200802",
x"E8B00003",
x"44A00006",
x"08002733",
x"44A00007",
x"E806005D",
x"44250803",
x"E8300003",
x"44200006",
x"08002739",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"0800273E",
x"2003FFFF",
x"08002740",
x"20030001",
x"48600003",
x"44002006",
x"08002744",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44611003",
x"47200802",
x"47421000",
x"44220803",
x"2004004C",
x"C4820000",
x"44401002",
x"47010800",
x"44410803",
x"46E10800",
x"44010003",
x"46200000",
x"44800003",
x"68030006",
x"68600003",
x"44000806",
x"08002789",
x"47E00801",
x"0800278B",
x"46C00801",
x"20030044",
x"C4600000",
x"44200002",
x"441E0003",
x"08002792",
x"20030088",
x"C4600000",
x"E4200008",
x"40210010",
x"C0000051",
x"20210010",
x"44000806",
x"C4200008",
x"44010001",
x"2003003C",
x"C4620000",
x"46A70801",
x"44210802",
x"44410801",
x"46A00001",
x"44000002",
x"44200801",
x"E8300003",
x"44200006",
x"080027A5",
x"46000006",
x"47600802",
x"20030038",
x"C4600000",
x"44200003",
x"E7E00230",
x"080027AB",
x"200C0000",
x"8FED0204",
x"40210010",
x"C0001777",
x"20210010",
x"48600025",
x"C7E1022C",
x"C7E00134",
x"44201002",
x"C7E10228",
x"C7E00130",
x"44200002",
x"44401000",
x"C7E10224",
x"C7E0012C",
x"44200002",
x"44400800",
x"44200807",
x"EA010003",
x"46000006",
x"080027C1",
x"44200006",
x"45400802",
x"8DC3FFE4",
x"C4600000",
x"44200002",
x"C7E20244",
x"C7E10238",
x"44010802",
x"44410800",
x"E7E10244",
x"C7E20240",
x"C7E10234",
x"44010802",
x"44410800",
x"E7E10240",
x"C7E2023C",
x"C7E10230",
x"44010002",
x"44400000",
x"E7E0023C",
x"E0000000",
x"E0000000",
x"6B200090",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"080027F8",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"43390002",
x"6B20006C",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"0800281B",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"43390002",
x"6B200048",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"0800283E",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"43390002",
x"6B200024",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"08002861",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C00024D7",
x"20210004",
x"43390002",
x"080027D6",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"20030004",
x"687A03E8",
x"A3430002",
x"4DA31800",
x"686003E4",
x"A3430002",
x"4D831800",
x"AC390000",
x"AC290004",
x"AC2A0008",
x"AC2B000C",
x"AC2C0010",
x"AC2D0014",
x"AC2E0018",
x"AC2F001C",
x"48600002",
x"08002C45",
x"A3430002",
x"4D431800",
x"C4600000",
x"E7E00244",
x"C460FFFC",
x"E7E00240",
x"C460FFF8",
x"E7E0023C",
x"8D3E0000",
x"A3430002",
x"4F23B000",
x"A3430002",
x"4DC3C000",
x"AC2B0020",
x"AC360024",
x"AC380028",
x"4BC00002",
x"08002941",
x"8FF702CC",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"080028DF",
x"20050002",
x"68A60002",
x"080028DF",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"080028D9",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"080028DE",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C00013F1",
x"20210030",
x"080028E5",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002902",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"0800291F",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"0800293C",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00027D6",
x"20210030",
x"4BDC0002",
x"080029FC",
x"8FF702C8",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08002999",
x"20050002",
x"68A60002",
x"08002999",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08002993",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08002998",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C00013F1",
x"20210030",
x"0800299F",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"080029BD",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"080029DA",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"080029F7",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00027D6",
x"20210030",
x"20030002",
x"4BC30002",
x"08002AB8",
x"8FF702C4",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08002A55",
x"20050002",
x"68A60002",
x"08002A55",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08002A4F",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08002A54",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C00013F1",
x"20210030",
x"08002A5B",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002A79",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002A96",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002AB3",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00027D6",
x"20210030",
x"20030003",
x"4BC30002",
x"08002B74",
x"8FF702C0",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08002B11",
x"20050002",
x"68A60002",
x"08002B11",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08002B0B",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08002B10",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C00013F1",
x"20210030",
x"08002B17",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002B35",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002B52",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002B6F",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00027D6",
x"20210030",
x"20030004",
x"4BC30002",
x"08002C30",
x"8FF702BC",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08002BCD",
x"20050002",
x"68A60002",
x"08002BCD",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08002BC7",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08002BCC",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C00013F1",
x"20210030",
x"08002BD3",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002BF1",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002C0E",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"08002C2B",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C00024D7",
x"20210030",
x"201E0070",
x"23D90000",
x"40210030",
x"C00027D6",
x"20210030",
x"A3430002",
x"8C2B0020",
x"4D631800",
x"C7E20250",
x"C4610000",
x"C7E00244",
x"44200002",
x"44400000",
x"E7E00250",
x"C7E2024C",
x"C461FFFC",
x"C7E00240",
x"44200002",
x"44400000",
x"E7E0024C",
x"C7E20248",
x"C461FFF8",
x"C7E0023C",
x"44200002",
x"44400000",
x"E7E00248",
x"235A0001",
x"8C2F001C",
x"8C2E0018",
x"8C2D0014",
x"8C2C0010",
x"8C2B000C",
x"8C2A0008",
x"8C290004",
x"8C390000",
x"08002867",
x"E0000000",
x"E0000000",
x"A0830002",
x"4CA33000",
x"20030004",
x"687A00A0",
x"8CC7FFF8",
x"A3430002",
x"4CE31800",
x"6860009B",
x"A0870002",
x"4D273800",
x"8CECFFF8",
x"A34B0002",
x"4D8B5800",
x"4963001D",
x"A08B0002",
x"4D0B5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"49630015",
x"408B0001",
x"A16B0002",
x"4CAB5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"4963000C",
x"208B0001",
x"A16B0002",
x"4CAB5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"49630003",
x"200B0001",
x"08002C76",
x"200B0000",
x"08002C78",
x"200B0000",
x"08002C7A",
x"200B0000",
x"08002C7C",
x"200B0000",
x"4960000C",
x"A0830002",
x"4CA31800",
x"8C79FFE4",
x"8C69FFE8",
x"8C6AFFEC",
x"8C6BFFF0",
x"8C6CFFF4",
x"8C6DFFF8",
x"8C6EFFFC",
x"8C6F0000",
x"08002867",
x"8CCBFFF4",
x"A3430002",
x"4D631800",
x"48600002",
x"08002CF1",
x"8CE7FFEC",
x"40830001",
x"A0630002",
x"4CA31800",
x"8C6BFFEC",
x"8CC6FFEC",
x"20830001",
x"A0630002",
x"4CA31800",
x"8C6CFFEC",
x"A0830002",
x"4D031800",
x"8C6DFFEC",
x"A3430002",
x"4CE31800",
x"C4600000",
x"E7E00244",
x"C460FFFC",
x"E7E00240",
x"C460FFF8",
x"E7E0023C",
x"A3430002",
x"4D631800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4CC31800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4D831800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4DA31800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A0830002",
x"4CA31800",
x"8C66FFF0",
x"A3430002",
x"4CC31800",
x"C7E20250",
x"C4610000",
x"C7E00244",
x"44200002",
x"44400000",
x"E7E00250",
x"C7E2024C",
x"C461FFFC",
x"C7E00240",
x"44200002",
x"44400000",
x"E7E0024C",
x"C7E20248",
x"C461FFF8",
x"C7E0023C",
x"44200002",
x"44400000",
x"E7E00248",
x"235A0001",
x"08002C51",
x"E0000000",
x"E0000000",
x"20030004",
x"687A00E2",
x"A3430002",
x"4D631800",
x"686000DE",
x"A3430002",
x"4D431800",
x"AC390000",
x"AC2D0004",
x"AC2A0008",
x"AC2B000C",
x"AC2C0010",
x"AC2E0014",
x"48600002",
x"08002DCF",
x"8F230000",
x"E7F00244",
x"E7F00240",
x"E7F0023C",
x"A0630002",
x"03E31820",
x"8C7702CC",
x"A3430002",
x"4FC3B000",
x"A3430002",
x"4D83C000",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40670001",
x"68E00052",
x"A0E30002",
x"03E31820",
x"8C630110",
x"8C66FFD8",
x"8C65FFFC",
x"C7010000",
x"8C64FFEC",
x"C4800000",
x"44200001",
x"E4C00000",
x"C701FFFC",
x"C480FFFC",
x"44200001",
x"E4C0FFFC",
x"C701FFF8",
x"C480FFF8",
x"44200001",
x"E4C0FFF8",
x"20040002",
x"48A4000F",
x"8C63FFF0",
x"C4C10000",
x"C4C3FFFC",
x"C4C2FFF8",
x"C4600000",
x"44010802",
x"C460FFFC",
x"44030002",
x"44200800",
x"C460FFF8",
x"44020002",
x"44200000",
x"E4C0FFF4",
x"08002D63",
x"20040002",
x"68850002",
x"08002D63",
x"C4C20000",
x"C4C1FFFC",
x"C4C0FFF8",
x"44422002",
x"8C64FFF0",
x"C4830000",
x"44832802",
x"44212002",
x"C483FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C483FFF8",
x"44831802",
x"44A32000",
x"8C64FFF4",
x"48800003",
x"44801806",
x"08002D5D",
x"44202802",
x"8C63FFDC",
x"C4630000",
x"44A31802",
x"44832000",
x"44021802",
x"C460FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C460FFF8",
x"44201802",
x"44831800",
x"20030003",
x"48A30003",
x"44710001",
x"08002D62",
x"44600006",
x"E4C0FFF4",
x"40E40001",
x"23030000",
x"4021001C",
x"C00013F1",
x"2021001C",
x"08002D69",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"AC290018",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"08002D87",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"08002DA4",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"08002DC1",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C00024D7",
x"20210020",
x"20030070",
x"20790000",
x"40210020",
x"C00027D6",
x"20210020",
x"8C290018",
x"A3430002",
x"4D231800",
x"C7E00244",
x"E4600000",
x"C7E00240",
x"E460FFFC",
x"C7E0023C",
x"E460FFF8",
x"235A0001",
x"8C2E0014",
x"8C2C0010",
x"8C2B000C",
x"8C2A0008",
x"8C2D0004",
x"8C390000",
x"08002CF5",
x"E0000000",
x"E0000000",
x"68C00076",
x"C7E30264",
x"8FE30260",
x"00C31822",
x"40210004",
x"C0000081",
x"20210004",
x"44600002",
x"C7E10288",
x"44010802",
x"442D0800",
x"E7E102AC",
x"C7E10284",
x"44010802",
x"442C0800",
x"E7E102A8",
x"C7E10280",
x"44010002",
x"440B0000",
x"E7E002A4",
x"C7E202AC",
x"44420802",
x"C7E002A8",
x"44000002",
x"44200800",
x"C7E002A4",
x"44000002",
x"44200000",
x"44000004",
x"C8100003",
x"46200803",
x"08002DFB",
x"200300C8",
x"C4610000",
x"44410002",
x"E7E002AC",
x"C7E002A8",
x"44010002",
x"E7E002A8",
x"C7E002A4",
x"44010002",
x"E7E002A4",
x"E7F00250",
x"E7F0024C",
x"E7F00248",
x"C7E00128",
x"E7E00270",
x"C7E00124",
x"E7E0026C",
x"C7E00120",
x"E7E00268",
x"20190000",
x"A0C30002",
x"4CE31800",
x"8C70FFE4",
x"8C75FFE8",
x"8C77FFEC",
x"8C71FFF0",
x"8C72FFF4",
x"8C73FFF8",
x"8C74FFFC",
x"8C780000",
x"43F602AC",
x"E42B0000",
x"E42C0004",
x"E42D0008",
x"AC28000C",
x"AC270010",
x"AC260014",
x"46007006",
x"46206806",
x"4021001C",
x"C00020C0",
x"2021001C",
x"8C260014",
x"A0C30002",
x"8C270010",
x"4CE31800",
x"8C630000",
x"C7E00250",
x"E4600000",
x"C7E0024C",
x"E460FFFC",
x"C7E00248",
x"E460FFF8",
x"A0C30002",
x"4CE31800",
x"8C63FFE8",
x"8C28000C",
x"AC680000",
x"A0C30002",
x"4CE31800",
x"201A0000",
x"8C7EFFE4",
x"8C79FFE8",
x"8C69FFEC",
x"8C6DFFF0",
x"8C6AFFF4",
x"8C6BFFF8",
x"8C6CFFFC",
x"8C6E0000",
x"4021001C",
x"C0002CF5",
x"2021001C",
x"8C260014",
x"40C60001",
x"8C28000C",
x"21030001",
x"20080005",
x"68680003",
x"40680005",
x"08002E4A",
x"20680000",
x"C42D0008",
x"C42C0004",
x"C42B0000",
x"8C270010",
x"08002DD9",
x"E0000000",
x"8FE30258",
x"68C30002",
x"E0000000",
x"A0C30002",
x"4CE31800",
x"8C630000",
x"C4600000",
x"E7E00250",
x"C460FFFC",
x"E7E0024C",
x"C460FFF8",
x"E7E00248",
x"8FE40254",
x"21430001",
x"68640003",
x"20030000",
x"08002E6D",
x"680A0003",
x"20030000",
x"08002E6D",
x"8FE40258",
x"20C30001",
x"68640003",
x"20030000",
x"08002E6D",
x"68060003",
x"20030000",
x"08002E6D",
x"20030001",
x"AC280000",
x"AC270004",
x"AC290008",
x"AC2A000C",
x"AC260010",
x"48600012",
x"A0C30002",
x"4CE32800",
x"201A0000",
x"8CB9FFE4",
x"8CA3FFE8",
x"8CA4FFEC",
x"8CABFFF0",
x"8CACFFF4",
x"8CADFFF8",
x"8CAEFFFC",
x"8CAF0000",
x"20690000",
x"208A0000",
x"40210018",
x"C0002867",
x"20210018",
x"08002E8A",
x"201A0000",
x"20E50000",
x"20C40000",
x"40210018",
x"C0002C51",
x"20210018",
x"C7E00250",
x"40210018",
x"C00000A0",
x"20210018",
x"20640000",
x"200300FF",
x"68640006",
x"68800003",
x"20830000",
x"08002E95",
x"20030000",
x"08002E97",
x"200300FF",
x"04600001",
x"C7E0024C",
x"40210018",
x"C00000A0",
x"20210018",
x"20640000",
x"200300FF",
x"68640006",
x"68800003",
x"20830000",
x"08002EA3",
x"20030000",
x"08002EA5",
x"200300FF",
x"04600001",
x"C7E00248",
x"40210018",
x"C00000A0",
x"20210018",
x"20640000",
x"200300FF",
x"68640006",
x"68800003",
x"20830000",
x"08002EB1",
x"20030000",
x"08002EB3",
x"200300FF",
x"04600001",
x"8C260010",
x"20C60001",
x"8C2A000C",
x"8C290008",
x"8C270004",
x"8C280000",
x"08002E50",
x"8FE40254",
x"69440002",
x"E0000000",
x"40840001",
x"AC230000",
x"AC280004",
x"AC290008",
x"AC27000C",
x"AC2A0010",
x"69440002",
x"08002EE3",
x"21450001",
x"C7E30264",
x"8FE4025C",
x"00A43022",
x"20C30000",
x"40210018",
x"C0000081",
x"20210018",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE40258",
x"40860001",
x"8C230000",
x"21070000",
x"20680000",
x"40210018",
x"C0002DD9",
x"20210018",
x"20060000",
x"8C2A0010",
x"8C27000C",
x"8C290008",
x"8C280004",
x"20FB0000",
x"21270000",
x"23690000",
x"40210018",
x"C0002E50",
x"20210018",
x"8C2A0010",
x"214A0001",
x"8C230000",
x"20630002",
x"20060005",
x"68660003",
x"40660005",
x"08002EF7",
x"20660000",
x"8FE30254",
x"69430002",
x"E0000000",
x"40630001",
x"AC260014",
x"AC2A0018",
x"69430002",
x"08002F1B",
x"21440001",
x"C7E30264",
x"8FE3025C",
x"00831822",
x"40210020",
x"C0000081",
x"20210020",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40630001",
x"8C27000C",
x"20C80000",
x"20660000",
x"40210020",
x"C0002DD9",
x"20210020",
x"20030000",
x"8C2A0018",
x"8C290008",
x"8C280004",
x"8C27000C",
x"20660000",
x"211B0000",
x"20E80000",
x"23670000",
x"40210020",
x"C0002E50",
x"20210020",
x"8C2A0018",
x"214A0001",
x"8C260014",
x"20C40002",
x"20030005",
x"68830003",
x"40830005",
x"08002F30",
x"20830000",
x"8C280004",
x"8C27000C",
x"8C290008",
x"211B0000",
x"21280000",
x"20E90000",
x"23670000",
x"08002EBB",
x"6920007D",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"206D0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20680000",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF0",
x"20030005",
x"20040000",
x"C000003F",
x"206C0000",
x"20030005",
x"20040000",
x"C000003F",
x"206B0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20670000",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF0",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20660000",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF0",
x"20030001",
x"20040000",
x"C000003F",
x"206E0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20650000",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"20210004",
x"ACA3FFF0",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6EFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC6BFFF4",
x"AC6CFFF8",
x"AC68FFFC",
x"AC6D0000",
x"A1240002",
x"6D441800",
x"41290001",
x"08002F38",
x"21430000",
x"E0000000",
x"E4200000",
x"E4220004",
x"20060005",
x"68860039",
x"44A51002",
x"44210002",
x"44400000",
x"44110000",
x"44000004",
x"44A01003",
x"44200803",
x"46200003",
x"A0A40002",
x"03E42020",
x"8C8502CC",
x"A0640002",
x"4CA42000",
x"8C840000",
x"E4820000",
x"E481FFFC",
x"E480FFF8",
x"20640028",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44202007",
x"E4820000",
x"E480FFFC",
x"E484FFF8",
x"20640050",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44401807",
x"E4800000",
x"E483FFFC",
x"E484FFF8",
x"20640001",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44000007",
x"E4830000",
x"E484FFFC",
x"E480FFF8",
x"20640029",
x"A0840002",
x"4CA42000",
x"8C840000",
x"E4830000",
x"E480FFFC",
x"E481FFF8",
x"20630051",
x"A0630002",
x"4CA31800",
x"8C630000",
x"E4600000",
x"E462FFFC",
x"E461FFF8",
x"E0000000",
x"44210002",
x"200600A4",
x"C4C60000",
x"44060000",
x"44002804",
x"46250003",
x"EA200006",
x"E8140003",
x"20060000",
x"08002FFE",
x"2006FFFF",
x"08003000",
x"20060001",
x"48C00003",
x"44002006",
x"08003004",
x"46202003",
x"44840002",
x"20070084",
x"C4EE0000",
x"45C00802",
x"20070080",
x"C4EF0000",
x"442F1803",
x"2007007C",
x"C4E10000",
x"E4210008",
x"C4210008",
x"44201002",
x"20070078",
x"C4E10000",
x"E421000C",
x"C421000C",
x"44230800",
x"44410803",
x"20070074",
x"C4EB0000",
x"45601002",
x"20070070",
x"C4ED0000",
x"45A10800",
x"44411003",
x"2007006C",
x"C4EC0000",
x"45801802",
x"20070068",
x"C4E10000",
x"E4210010",
x"C4210010",
x"44220800",
x"44610803",
x"20070064",
x"C4E90000",
x"45201002",
x"47810800",
x"44411003",
x"20070060",
x"C4EA0000",
x"45401802",
x"2007005C",
x"C4E10000",
x"E4210014",
x"C4210014",
x"44220800",
x"44611003",
x"2007004C",
x"C4E10000",
x"E4210018",
x"20070058",
x"C4E80000",
x"45001802",
x"20070054",
x"C4E10000",
x"E421001C",
x"C421001C",
x"44220800",
x"44610803",
x"20070050",
x"C4E70000",
x"44E01002",
x"47210800",
x"44410803",
x"47201002",
x"47410800",
x"44411003",
x"C4210018",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800803",
x"68060006",
x"68C00003",
x"44200006",
x"08003055",
x"47E10001",
x"08003057",
x"46C10001",
x"C4210004",
x"44010802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44052802",
x"20840001",
x"44A50002",
x"44060000",
x"44003004",
x"46260003",
x"EA200006",
x"E8140003",
x"20060000",
x"0800306E",
x"2006FFFF",
x"08003070",
x"20060001",
x"48C00003",
x"44000806",
x"08003074",
x"46200803",
x"44210002",
x"45C01002",
x"444F1803",
x"C4220008",
x"44402002",
x"C422000C",
x"44431000",
x"44821003",
x"45601802",
x"45A21000",
x"44621803",
x"45802002",
x"C4220010",
x"44431000",
x"44821003",
x"45201802",
x"47821000",
x"44621003",
x"45401802",
x"C4240014",
x"44821000",
x"44621003",
x"45002002",
x"C423001C",
x"44621000",
x"44821003",
x"44E01802",
x"47221000",
x"44621003",
x"47201802",
x"47421000",
x"44621003",
x"C4230018",
x"44601802",
x"47021000",
x"44621003",
x"46E21000",
x"44020003",
x"46200000",
x"44200803",
x"68060006",
x"68C00003",
x"44200006",
x"080030A1",
x"47E10001",
x"080030A3",
x"46C10001",
x"C4210000",
x"44010002",
x"44001002",
x"44590803",
x"47410801",
x"44410803",
x"47010801",
x"44410803",
x"46E10801",
x"44410803",
x"46210801",
x"44010003",
x"44060802",
x"C4220004",
x"C4200000",
x"08002FB7",
x"694000AA",
x"E4200000",
x"21430000",
x"40210008",
x"C0000081",
x"20210008",
x"44000806",
x"200300AC",
x"C4650000",
x"44250802",
x"200300A8",
x"C4640000",
x"44241001",
x"20040000",
x"C4200000",
x"E4240004",
x"E4250008",
x"E421000C",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210014",
x"C0002FB7",
x"20210014",
x"200300A4",
x"C4630000",
x"C421000C",
x"44231000",
x"20040000",
x"210B0002",
x"C4200000",
x"E4230010",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210018",
x"C0002FB7",
x"20210018",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"080030E2",
x"20690000",
x"6940007A",
x"21430000",
x"40210018",
x"C0000081",
x"20210018",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E4210014",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"4021001C",
x"C0002FB7",
x"2021001C",
x"C4230010",
x"C4210014",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"4021001C",
x"C0002FB7",
x"2021001C",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003109",
x"20690000",
x"69400052",
x"21430000",
x"4021001C",
x"C0000081",
x"2021001C",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E4210018",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210020",
x"C0002FB7",
x"20210020",
x"C4230010",
x"C4210018",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210020",
x"C0002FB7",
x"20210020",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003130",
x"20690000",
x"6940002A",
x"21430000",
x"40210020",
x"C0000081",
x"20210020",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E421001C",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210024",
x"C0002FB7",
x"20210024",
x"C4230010",
x"C421001C",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210024",
x"C0002FB7",
x"20210024",
x"414A0001",
x"21240001",
x"20030005",
x"68830003",
x"40830005",
x"08003157",
x"20830000",
x"C4200000",
x"20690000",
x"080030B3",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"69A00132",
x"21A30000",
x"40210004",
x"C0000081",
x"20210004",
x"200300AC",
x"C4640000",
x"44040002",
x"200300A8",
x"C4630000",
x"44030001",
x"20030004",
x"E4200000",
x"40210008",
x"C0000081",
x"20210008",
x"44000806",
x"44240802",
x"44235001",
x"20040000",
x"C4200000",
x"E42A0004",
x"E4230008",
x"E424000C",
x"E4210010",
x"21030000",
x"21850000",
x"45401006",
x"46000806",
x"46002806",
x"40210018",
x"C0002FB7",
x"20210018",
x"200300A4",
x"C4650000",
x"C4210010",
x"44254800",
x"20040000",
x"210A0002",
x"C4200000",
x"E4290014",
x"E4250018",
x"21430000",
x"21850000",
x"45201006",
x"46000806",
x"46002806",
x"40210020",
x"C0002FB7",
x"20210020",
x"20060003",
x"21830001",
x"20090005",
x"68690003",
x"40690005",
x"08003197",
x"20690000",
x"20C30000",
x"40210020",
x"C0000081",
x"20210020",
x"44000806",
x"C424000C",
x"44240802",
x"C4230008",
x"44234001",
x"20040000",
x"C4200000",
x"E428001C",
x"E4210020",
x"21030000",
x"21250000",
x"45001006",
x"46000806",
x"46002806",
x"40210028",
x"C0002FB7",
x"20210028",
x"C4250018",
x"C4210020",
x"44253800",
x"20040000",
x"C4200000",
x"E4270024",
x"21430000",
x"21250000",
x"44E01006",
x"46000806",
x"46002806",
x"4021002C",
x"C0002FB7",
x"2021002C",
x"20060002",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"080031C1",
x"20690000",
x"20C30000",
x"4021002C",
x"C0000081",
x"2021002C",
x"44000806",
x"C424000C",
x"44240802",
x"C4230008",
x"44233001",
x"20040000",
x"C4200000",
x"E4260028",
x"E421002C",
x"21030000",
x"21250000",
x"44C01006",
x"46000806",
x"46002806",
x"40210034",
x"C0002FB7",
x"20210034",
x"C4250018",
x"C421002C",
x"44251000",
x"20040000",
x"C4200000",
x"E4220030",
x"21430000",
x"21250000",
x"46000806",
x"46002806",
x"40210038",
x"C0002FB7",
x"20210038",
x"20060001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"080031EA",
x"20690000",
x"20C30000",
x"40210038",
x"C0000081",
x"20210038",
x"44000806",
x"C424000C",
x"44245802",
x"C4230008",
x"45630801",
x"20040000",
x"C4200000",
x"E42B0034",
x"21030000",
x"21250000",
x"44201006",
x"46002806",
x"46000806",
x"4021003C",
x"C0002FB7",
x"2021003C",
x"C4250018",
x"C42B0034",
x"45650800",
x"20040000",
x"C4200000",
x"21430000",
x"21250000",
x"44201006",
x"46002806",
x"46000806",
x"4021003C",
x"C0002FB7",
x"2021003C",
x"200A0000",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003212",
x"20690000",
x"C4200000",
x"AC280038",
x"40210040",
x"C00030B3",
x"20210040",
x"41AE0001",
x"21830002",
x"200C0005",
x"686C0003",
x"406C0005",
x"0800321E",
x"206C0000",
x"8C280038",
x"210D0004",
x"69C0006F",
x"21C30000",
x"40210040",
x"C0000081",
x"20210040",
x"C424000C",
x"44040002",
x"C4230008",
x"44030001",
x"20040000",
x"C42A0004",
x"E420003C",
x"21A30000",
x"21850000",
x"45401006",
x"46000806",
x"46002806",
x"40210044",
x"C0002FB7",
x"20210044",
x"20040000",
x"21A80002",
x"C4290014",
x"C420003C",
x"21030000",
x"21850000",
x"45201006",
x"46000806",
x"46002806",
x"40210044",
x"C0002FB7",
x"20210044",
x"21830001",
x"20050005",
x"68650003",
x"40650005",
x"08003246",
x"20650000",
x"20040000",
x"C428001C",
x"C420003C",
x"AC250040",
x"21A30000",
x"45001006",
x"46000806",
x"46002806",
x"40210048",
x"C0002FB7",
x"20210048",
x"20040000",
x"C4270024",
x"C420003C",
x"8C250040",
x"21030000",
x"44E01006",
x"46000806",
x"46002806",
x"40210048",
x"C0002FB7",
x"20210048",
x"8C250040",
x"20A30001",
x"20050005",
x"68650003",
x"40650005",
x"08003263",
x"20650000",
x"20040000",
x"C4260028",
x"C420003C",
x"AC250044",
x"21A30000",
x"44C01006",
x"46000806",
x"46002806",
x"4021004C",
x"C0002FB7",
x"2021004C",
x"20040000",
x"C4220030",
x"C420003C",
x"8C250044",
x"21030000",
x"46000806",
x"46002806",
x"4021004C",
x"C0002FB7",
x"2021004C",
x"200A0001",
x"8C250044",
x"20A30001",
x"20090005",
x"68690003",
x"40690005",
x"08003280",
x"20690000",
x"C420003C",
x"21A80000",
x"4021004C",
x"C00030B3",
x"2021004C",
x"41C40001",
x"21830002",
x"200C0005",
x"686C0003",
x"406C0005",
x"0800328C",
x"206C0000",
x"21A80004",
x"208D0000",
x"0800315E",
x"E0000000",
x"E0000000",
x"68E00058",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20640000",
x"8FE3001C",
x"AC240000",
x"40210008",
x"C000003F",
x"20210008",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240000",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E00042",
x"20030003",
x"46000006",
x"40210008",
x"C0000048",
x"20210008",
x"20640000",
x"8FE3001C",
x"AC240004",
x"4021000C",
x"C000003F",
x"2021000C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240004",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E0002C",
x"20030003",
x"46000006",
x"4021000C",
x"C0000048",
x"2021000C",
x"20640000",
x"8FE3001C",
x"AC240008",
x"40210010",
x"C000003F",
x"20210010",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240008",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E00016",
x"20030003",
x"46000006",
x"40210010",
x"C0000048",
x"20210010",
x"20640000",
x"8FE3001C",
x"AC24000C",
x"40210014",
x"C000003F",
x"20210014",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24000C",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"08003291",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"690000C2",
x"20060078",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20640000",
x"8FE3001C",
x"AC240000",
x"40210008",
x"C000003F",
x"20210008",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240000",
x"AC640000",
x"20640000",
x"20C30000",
x"40210008",
x"C000003F",
x"A1040002",
x"03E42020",
x"AC8302CC",
x"A1030002",
x"03E31820",
x"8C6602CC",
x"20030003",
x"46000006",
x"C0000048",
x"20210008",
x"20640000",
x"8FE3001C",
x"AC240004",
x"4021000C",
x"C000003F",
x"2021000C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240004",
x"AC640000",
x"ACC3FE28",
x"20030003",
x"46000006",
x"4021000C",
x"C0000048",
x"2021000C",
x"20640000",
x"8FE3001C",
x"AC240008",
x"40210010",
x"C000003F",
x"20210010",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240008",
x"AC640000",
x"ACC3FE2C",
x"20030003",
x"46000006",
x"40210010",
x"C0000048",
x"20210010",
x"20640000",
x"8FE3001C",
x"AC24000C",
x"40210014",
x"C000003F",
x"20210014",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24000C",
x"AC640000",
x"ACC3FE30",
x"20030003",
x"46000006",
x"40210014",
x"C0000048",
x"20210014",
x"20640000",
x"8FE3001C",
x"AC240010",
x"40210018",
x"C000003F",
x"20210018",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240010",
x"AC640000",
x"ACC3FE34",
x"20070072",
x"40210018",
x"C0003291",
x"20210018",
x"41080001",
x"69000058",
x"20060078",
x"20030003",
x"46000006",
x"40210018",
x"C0000048",
x"20210018",
x"20640000",
x"8FE3001C",
x"AC240014",
x"4021001C",
x"C000003F",
x"2021001C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240014",
x"AC640000",
x"20640000",
x"20C30000",
x"4021001C",
x"C000003F",
x"A1040002",
x"03E42020",
x"AC8302CC",
x"A1030002",
x"03E31820",
x"8C6602CC",
x"20030003",
x"46000006",
x"C0000048",
x"2021001C",
x"20640000",
x"8FE3001C",
x"AC240018",
x"40210020",
x"C000003F",
x"20210020",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240018",
x"AC640000",
x"ACC3FE28",
x"20030003",
x"46000006",
x"40210020",
x"C0000048",
x"20210020",
x"20640000",
x"8FE3001C",
x"AC24001C",
x"40210024",
x"C000003F",
x"20210024",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24001C",
x"AC640000",
x"ACC3FE2C",
x"20030003",
x"46000006",
x"40210024",
x"C0000048",
x"20210024",
x"20640000",
x"8FE3001C",
x"AC240020",
x"40210028",
x"C000003F",
x"20210028",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240020",
x"AC640000",
x"ACC3FE30",
x"20070073",
x"40210028",
x"C0003291",
x"20210028",
x"41080001",
x"080032EA",
x"E0000000",
x"E0000000",
x"69800060",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"69800054",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"69800048",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"6980003C",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"69800030",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"69800024",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"69800018",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"6980000C",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"20210004",
x"418C0001",
x"080033AD",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"69A0006E",
x"A1A30002",
x"03E31820",
x"8C6B02CC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE40",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"200C006F",
x"C00033AD",
x"20210004",
x"41AD0001",
x"69A00034",
x"A1A30002",
x"03E31820",
x"8C6B02CC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C000132A",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C000132A",
x"200C0070",
x"C00033AD",
x"20210004",
x"41AD0001",
x"0800340E",
x"E0000000",
x"E0000000",
x"00000000"

	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



