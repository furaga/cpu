library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is
	port (
		clka : in std_logic;
		addra : in std_logic_vector(13 downto 0);
		douta : out std_logic_vector(31 downto 0));



end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 1023) of word_t;
	signal addr_in	: integer range 0 to 1023;

	constant mem : mem_t := (
x"000000F4",
x"00000000",
x"3F800000",
x"BF800000",
x"00800000",
x"4B000000",
x"4B000000",
x"43160000",
x"C3160000",
x"C0000000",
x"3B800000",
x"41A00000",
x"3D4CCCC4",
x"3E800000",
x"41200000",
x"3E999999",
x"3E199999",
x"40490FDA",
x"41F00000",
x"BFC90FDA",
x"40800000",
x"41800000",
x"41300000",
x"41C80000",
x"41500000",
x"42100000",
x"42440000",
x"41880000",
x"42800000",
x"41980000",
x"42A20000",
x"41A80000",
x"42C80000",
x"41B80000",
x"42F20000",
x"41700000",
x"38D1B70F",
x"4CBEBC20",
x"BDCCCCC4",
x"3C23D70A",
x"BE4CCCC4",
x"BF800000",
x"3DCCCCC4",
x"3F66665E",
x"3E4CCCC4",
x"C3480000",
x"43480000",
x"40400000",
x"40A00000",
x"41100000",
x"40E00000",
x"3F800000",
x"3C8EFA2D",
x"43000000",
x"4E6E6B28",
x"437F0000",
x"00000000",
x"3FC90FDA",
x"3F000000",
x"40C90FDA",
x"40000000",
x"40490FDA",
x"080000C2",
x"A0630002",
x"00622820",
x"20430000",
x"68A20005",
x"28A20004",
x"AC440000",
x"20420004",
x"08000042",
x"E0000000",
x"A0630002",
x"00622020",
x"20430000",
x"68820005",
x"28820004",
x"E4400000",
x"20420004",
x"0800004B",
x"E0000000",
x"44000806",
x"20030000",
x"C4640000",
x"E8800015",
x"C8800014",
x"44000007",
x"20030010",
x"C4620000",
x"E8020004",
x"C8020003",
x"44000007",
x"E0000000",
x"44020000",
x"44020001",
x"44200807",
x"E820001B",
x"C820001A",
x"44020000",
x"20030004",
x"C4630000",
x"44030000",
x"44020001",
x"44000007",
x"E0000000",
x"20030010",
x"C4620000",
x"E8020003",
x"C8020002",
x"E0000000",
x"44000806",
x"44020000",
x"E4200000",
x"8C240000",
x"44020001",
x"E4200000",
x"8C240000",
x"E8010005",
x"C8010004",
x"20030004",
x"C4630000",
x"44030001",
x"E0000000",
x"44000007",
x"E0000000",
x"44000007",
x"C0000051",
x"44000007",
x"E0000000",
x"68030006",
x"28030005",
x"00031822",
x"C0000087",
x"44000007",
x"E0000000",
x"20050010",
x"C4A10000",
x"20050014",
x"8CA40000",
x"2005000C",
x"8CA50000",
x"68A30007",
x"28A30006",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"E0000000",
x"20040000",
x"C4820000",
x"00651822",
x"44411000",
x"68A3FFFE",
x"28A3FFFD",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"44020000",
x"E0000000",
x"20030000",
x"C4610000",
x"E8200006",
x"C8200005",
x"44000007",
x"C00000A8",
x"00031822",
x"E0000000",
x"C0000051",
x"20040010",
x"C4820000",
x"20040014",
x"8C840000",
x"E8400007",
x"C8400006",
x"44020000",
x"E4200000",
x"8C230000",
x"00641822",
x"E0000000",
x"2005000C",
x"8CA50000",
x"20030000",
x"44020001",
x"00651820",
x"E840FFFE",
x"C840FFFD",
x"44020000",
x"E4200000",
x"8C250000",
x"00A42822",
x"00A31820",
x"E0000000",
x"080000A0",
x"203F0000",
x"40210948",
x"201C0001",
x"201DFFFF",
x"201B00DC",
x"C7700000",
x"201B00C8",
x"C7710000",
x"201B0018",
x"C7720000",
x"201B001C",
x"C7730000",
x"201B00A0",
x"C7740000",
x"201B00E4",
x"C7750000",
x"201B00E0",
x"C7760000",
x"201B00B8",
x"C7770000",
x"201B00BC",
x"C7780000",
x"201B00C0",
x"C7790000",
x"201B00C4",
x"C77A0000",
x"201B00D8",
x"C77B0000",
x"201B0088",
x"C77C0000",
x"201B00E8",
x"C77D0000",
x"201B0040",
x"C77E0000",
x"201B0048",
x"C77F0000",
x"200300F0",
x"C4650000",
x"200300EC",
x"C46A0000",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20004",
x"40210004",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20008",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E2000C",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20010",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040001",
x"AFE20944",
x"43E20014",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20018",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E2001C",
x"C000003F",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E20020",
x"46000006",
x"C0000048",
x"20640000",
x"8FE20944",
x"2006003C",
x"200A0000",
x"20090000",
x"20080000",
x"20070000",
x"20050000",
x"20430000",
x"2042002C",
x"AC64FFD8",
x"AC64FFDC",
x"AC64FFE0",
x"AC64FFE4",
x"AC65FFE8",
x"AC64FFEC",
x"AC64FFF0",
x"AC67FFF4",
x"AC68FFF8",
x"AC69FFFC",
x"AC6A0000",
x"AFE20944",
x"43E20110",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2011C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20128",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20134",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030001",
x"AFE20944",
x"43E20138",
x"47600006",
x"C0000048",
x"8FE20944",
x"20060032",
x"20030001",
x"2004FFFF",
x"C000003F",
x"20640000",
x"AFE20944",
x"43E20200",
x"20C30000",
x"C000003F",
x"8FE20944",
x"20060001",
x"20030001",
x"8FE40200",
x"C000003F",
x"20640000",
x"AFE20944",
x"43E20204",
x"20C30000",
x"C000003F",
x"8FE20944",
x"20030001",
x"AFE20944",
x"43E20208",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E2020C",
x"C000003F",
x"8FE20944",
x"20030001",
x"200400D4",
x"C4800000",
x"AFE20944",
x"43E20210",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2021C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20220",
x"C000003F",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2022C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20238",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20244",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20250",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030002",
x"20040000",
x"AFE20944",
x"43E20258",
x"C000003F",
x"8FE20944",
x"20030002",
x"20040000",
x"AFE20944",
x"43E20260",
x"C000003F",
x"8FE20944",
x"20030001",
x"AFE20944",
x"43E20264",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20270",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2027C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20288",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20294",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E202A0",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E202AC",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E202B0",
x"46000006",
x"C0000048",
x"20670000",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E202B4",
x"43E402B0",
x"C000003F",
x"20640000",
x"8FE20944",
x"20060000",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"AFE20944",
x"43E202B8",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E202CC",
x"43E402B8",
x"C000003F",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E202D0",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E202DC",
x"46000006",
x"C0000048",
x"20660000",
x"8FE20944",
x"2003003C",
x"AFE20944",
x"43E203CC",
x"43E402D0",
x"C000003F",
x"20640000",
x"8FE20944",
x"AFE20944",
x"43E203D4",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC660000",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E203D8",
x"46000006",
x"C0000048",
x"20660000",
x"8FE20944",
x"20030000",
x"AFE20944",
x"43E203DC",
x"43E403D8",
x"C000003F",
x"8FE20944",
x"AFE20944",
x"43E203E4",
x"20440000",
x"20420008",
x"AC83FFFC",
x"AC860000",
x"8FE20944",
x"200600B4",
x"20050000",
x"20430000",
x"2042000C",
x"E470FFF8",
x"AC64FFFC",
x"AC650000",
x"AFE20944",
x"43E206B4",
x"20640000",
x"20C30000",
x"C000003F",
x"8FE20944",
x"20030001",
x"20040000",
x"AFE20944",
x"43E206B8",
x"C000003F",
x"8FE20944",
x"20030080",
x"20040080",
x"AFE30258",
x"AFE40254",
x"20040040",
x"AFE40260",
x"20040040",
x"AFE4025C",
x"200400D0",
x"C4830000",
x"C0000081",
x"44600003",
x"E7E00264",
x"8FEC0258",
x"20030003",
x"AFE20944",
x"43E206C4",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E206D0",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E206E4",
x"43E406D0",
x"C000003F",
x"206A0000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306E0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306DC",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306D8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE306D4",
x"20030005",
x"20040000",
x"AFE20944",
x"43E206F8",
x"C000003F",
x"20690000",
x"8FE20944",
x"20030005",
x"20040000",
x"AFE20944",
x"43E2070C",
x"C000003F",
x"20680000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20718",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E2072C",
x"43E40718",
x"C000003F",
x"20670000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30728",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30724",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30720",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3071C",
x"20030003",
x"AFE20944",
x"43E20738",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E2074C",
x"43E40738",
x"C000003F",
x"20660000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30748",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30744",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30740",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3073C",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20750",
x"C000003F",
x"206D0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2075C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E20770",
x"43E4075C",
x"C000003F",
x"20650000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3076C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30768",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30764",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30760",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA0774",
x"8FE30258",
x"40690002",
x"C0003922",
x"20720000",
x"AFF20778",
x"8FEC0258",
x"20030003",
x"AFE20944",
x"43E20784",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20790",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E207A4",
x"43E40790",
x"C000003F",
x"206A0000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307A0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3079C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30798",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30794",
x"20030005",
x"20040000",
x"AFE20944",
x"43E207B8",
x"C000003F",
x"20690000",
x"8FE20944",
x"20030005",
x"20040000",
x"AFE20944",
x"43E207CC",
x"C000003F",
x"20680000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E207D8",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E207EC",
x"43E407D8",
x"C000003F",
x"20670000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307E0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307DC",
x"20030003",
x"AFE20944",
x"43E207F8",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E2080C",
x"43E407F8",
x"C000003F",
x"20660000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30808",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30804",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30800",
x"20030003",
x"46000006",
x"C0000048",
x"AFE307FC",
x"20030001",
x"20040000",
x"AFE20944",
x"43E20810",
x"C000003F",
x"206D0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E2081C",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E20830",
x"43E4081C",
x"C000003F",
x"20650000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3082C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30828",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30824",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30820",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA0834",
x"8FE30258",
x"40690002",
x"C0003922",
x"20700000",
x"AFF00838",
x"8FEC0258",
x"20030003",
x"AFE20944",
x"43E20844",
x"46000006",
x"C0000048",
x"206B0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20850",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E20864",
x"43E40850",
x"C000003F",
x"206A0000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30860",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3085C",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30858",
x"20030003",
x"46000006",
x"C0000048",
x"AFE30854",
x"20030005",
x"20040000",
x"AFE20944",
x"43E20878",
x"C000003F",
x"20690000",
x"8FE20944",
x"20030005",
x"20040000",
x"AFE20944",
x"43E2088C",
x"C000003F",
x"20680000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E20898",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E208AC",
x"43E40898",
x"C000003F",
x"20670000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308A0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE3089C",
x"20030003",
x"AFE20944",
x"43E208B8",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E208CC",
x"43E408B8",
x"C000003F",
x"20660000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308C0",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308BC",
x"20030001",
x"20040000",
x"AFE20944",
x"43E208D0",
x"C000003F",
x"206D0000",
x"8FE20944",
x"20030003",
x"AFE20944",
x"43E208DC",
x"46000006",
x"C0000048",
x"8FE20944",
x"20030005",
x"AFE20944",
x"43E208F0",
x"43E408DC",
x"C000003F",
x"20650000",
x"8FE20944",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308EC",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E8",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E4",
x"20030003",
x"46000006",
x"C0000048",
x"AFE308E0",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6DFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC68FFF4",
x"AC69FFF8",
x"AC6AFFFC",
x"AC6B0000",
x"20640000",
x"21830000",
x"C000003F",
x"206A0000",
x"AFEA08F4",
x"8FE30258",
x"40690002",
x"C0003922",
x"20210004",
x"20710000",
x"AFF108F8",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800043C",
x"20030001",
x"0800043E",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08000444",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08000454",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800045E",
x"20040001",
x"08000460",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08000476",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08000487",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800048C",
x"44000807",
x"E7E1011C",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800049D",
x"20030001",
x"0800049F",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080004A5",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080004B5",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080004BF",
x"20040001",
x"080004C1",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080004D7",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"080004E8",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080004ED",
x"44000807",
x"E7E10118",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080004FE",
x"20030001",
x"08000500",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08000506",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08000516",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000520",
x"20040001",
x"08000522",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08000538",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08000549",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800054E",
x"44000807",
x"E7E10114",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800055F",
x"20030001",
x"08000561",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08000567",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08000577",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000581",
x"20040001",
x"08000583",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08000599",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"080005AA",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080005AF",
x"44000807",
x"200300CC",
x"C4680000",
x"44281802",
x"46C31001",
x"E8500003",
x"44400806",
x"080005B7",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080005DD",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080005CE",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005C9",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080005CE",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080005DD",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005D8",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080005DD",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000600",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080005F1",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005EC",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080005F1",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000600",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080005FB",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000600",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA020003",
x"20030000",
x"08000605",
x"20030001",
x"0800060A",
x"EA020003",
x"20030001",
x"0800060A",
x"20030000",
x"E8A00003",
x"44000806",
x"0800060E",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000612",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44003807",
x"08000625",
x"44003806",
x"E8700003",
x"44600806",
x"08000629",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"0800064F",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000640",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800063B",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000640",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"0800064F",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800064A",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"0800064F",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000672",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000663",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800065E",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000663",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000672",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800066D",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000672",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA030003",
x"20030000",
x"08000677",
x"20030001",
x"0800067C",
x"EA030003",
x"20030001",
x"0800067C",
x"20030000",
x"E8A00003",
x"44000806",
x"08000680",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000684",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44003007",
x"08000697",
x"44003006",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080006A7",
x"20030001",
x"080006A9",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080006AF",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080006BF",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080006C9",
x"20040001",
x"080006CB",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080006E1",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"080006F2",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080006F7",
x"44000807",
x"44281802",
x"46C31001",
x"E8500003",
x"44400806",
x"080006FD",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000723",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000714",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800070F",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000714",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000723",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800071E",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000723",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000746",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000737",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000732",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000737",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000746",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000741",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000746",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA020003",
x"20030000",
x"0800074B",
x"20030001",
x"08000750",
x"EA020003",
x"20030001",
x"08000750",
x"20030000",
x"E8A00003",
x"44000806",
x"08000754",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000758",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44001007",
x"0800076B",
x"44001006",
x"E8700003",
x"44600806",
x"0800076F",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000795",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000786",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000781",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000786",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000795",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000790",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000795",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080007B8",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080007A9",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007A4",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080007A9",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080007B8",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080007B3",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080007B8",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA030003",
x"20030000",
x"080007BD",
x"20030001",
x"080007C2",
x"EA030003",
x"20030001",
x"080007C2",
x"20030000",
x"E8A00003",
x"44000806",
x"080007C6",
x"47A00801",
x"EAC10003",
x"44200006",
x"080007CA",
x"44A10001",
x"44150802",
x"44210002",
x"44191803",
x"47431801",
x"44031803",
x"47031801",
x"44031803",
x"46E31801",
x"44030003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"080007DD",
x"44200006",
x"44E01802",
x"200300B4",
x"C4610000",
x"44611802",
x"E7E302A0",
x"200300B0",
x"C4630000",
x"44C31802",
x"E7E3029C",
x"44E21802",
x"44610802",
x"E7E10298",
x"E7E20288",
x"E7F00284",
x"44000807",
x"E7E10280",
x"44C00807",
x"44200002",
x"E7E00294",
x"44E03807",
x"E7E70290",
x"44220002",
x"E7E0028C",
x"C7E1011C",
x"C7E002A0",
x"44200001",
x"E7E00128",
x"C7E10118",
x"C7E0029C",
x"44200001",
x"E7E00124",
x"C7E10114",
x"C7E00298",
x"44200001",
x"E7E00120",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800080C",
x"20030001",
x"0800080E",
x"20030001",
x"48600012",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08000814",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"08000824",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000834",
x"20030001",
x"08000836",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"0800083C",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"0800084C",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000856",
x"20040001",
x"08000858",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"0800086E",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"0800087F",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08000884",
x"44000807",
x"44281802",
x"E8700003",
x"44600806",
x"08000889",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080008AF",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080008A0",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800089B",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008A0",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008AF",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080008AA",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008AF",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008D2",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080008C3",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080008BE",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008C3",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008D2",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080008CD",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080008D2",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA030003",
x"20030000",
x"080008D7",
x"20030001",
x"080008DC",
x"EA030003",
x"20030001",
x"080008DC",
x"20030000",
x"E8A00003",
x"44000806",
x"080008E0",
x"47A00801",
x"EAC10003",
x"44200006",
x"080008E4",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"080008F7",
x"44200006",
x"44000007",
x"E7E00130",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000909",
x"20030001",
x"0800090B",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08000911",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08000921",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800092B",
x"20040001",
x"0800092D",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08000943",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44003006",
x"8FE30010",
x"C0000081",
x"44002006",
x"8FE30014",
x"C0000081",
x"20210004",
x"44800003",
x"44C00000",
x"08000954",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08000959",
x"44000807",
x"44282002",
x"46C31001",
x"E8500003",
x"44400806",
x"0800095F",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000985",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000976",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000971",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000976",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000985",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000980",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000985",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009A8",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000999",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000994",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000999",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009A8",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080009A3",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009A8",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA020003",
x"20030000",
x"080009AD",
x"20030001",
x"080009B2",
x"EA020003",
x"20030001",
x"080009B2",
x"20030000",
x"E8A00003",
x"44000806",
x"080009B6",
x"47A00801",
x"EAC10003",
x"44200006",
x"080009BA",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44001807",
x"080009CD",
x"44001806",
x"E8900003",
x"44800806",
x"080009D1",
x"44800807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080009F7",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080009E8",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080009E3",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009E8",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009F7",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080009F2",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"080009F7",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A1A",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000A0B",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A06",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A0B",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A1A",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A15",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A1A",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA040003",
x"20030000",
x"08000A1F",
x"20030001",
x"08000A24",
x"EA040003",
x"20030001",
x"08000A24",
x"20030000",
x"E8A00003",
x"44000806",
x"08000A28",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000A2C",
x"44A10001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"08000A3F",
x"44200006",
x"44600002",
x"E7E00134",
x"46C41001",
x"E8500003",
x"44400806",
x"08000A46",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08000A6C",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000A5D",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A58",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A5D",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A6C",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A67",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A6C",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A8F",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08000A80",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A7B",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A80",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A8F",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08000A8A",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08000A8F",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8A00006",
x"EA020003",
x"20030000",
x"08000A94",
x"20030001",
x"08000A99",
x"EA020003",
x"20030001",
x"08000A99",
x"20030000",
x"E8A00003",
x"44000806",
x"08000A9D",
x"47A00801",
x"EAC10003",
x"44200006",
x"08000AA1",
x"44A10001",
x"44150002",
x"44001002",
x"44590803",
x"47410801",
x"44410803",
x"47010801",
x"44410803",
x"46E10801",
x"44410803",
x"46210801",
x"44010003",
x"45400802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"08000AB4",
x"44200006",
x"44600002",
x"E7E0012C",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000AC6",
x"20030001",
x"08000AC8",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08000ACE",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08000ADE",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000AE8",
x"20040001",
x"08000AEA",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08000B00",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08000B11",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08000B16",
x"44000807",
x"E7E10138",
x"20130000",
x"AC300000",
x"E42A0004",
x"22700000",
x"4021000C",
x"C000110D",
x"2021000C",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200A0030",
x"68AA0007",
x"200A0039",
x"69450003",
x"200A0000",
x"08000B2A",
x"200A0001",
x"08000B2C",
x"200A0001",
x"49400013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08000B32",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"206A0000",
x"08000B44",
x"20060000",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"206A0000",
x"495D0007",
x"20030001",
x"2004FFFF",
x"4021000C",
x"C000003F",
x"2021000C",
x"08000B50",
x"20080001",
x"4021000C",
x"C0001AF7",
x"2021000C",
x"AC6A0000",
x"AFE308FC",
x"8C640000",
x"489D0002",
x"08000B59",
x"AFE30200",
x"200B0001",
x"4021000C",
x"C0001C2F",
x"2021000C",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000B65",
x"20030001",
x"08000B67",
x"20030001",
x"48600012",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08000B6D",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"08000B7D",
x"20060000",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"487D0008",
x"20030001",
x"2004FFFF",
x"4021000C",
x"C000003F",
x"2021000C",
x"20640000",
x"08000B8D",
x"20080001",
x"AC230008",
x"40210010",
x"C0001AF7",
x"20210010",
x"20640000",
x"8C230008",
x"AC830000",
x"AFE40900",
x"8C830000",
x"487D0006",
x"20030001",
x"40210010",
x"C000003F",
x"20210010",
x"08000B9C",
x"200B0001",
x"AC24000C",
x"40210014",
x"C0001BA6",
x"20210014",
x"8C24000C",
x"AC640000",
x"AFE30204",
x"20030050",
x"04600001",
x"20030033",
x"04600001",
x"2003000A",
x"04600001",
x"8FE40258",
x"40210014",
x"C0001037",
x"20030020",
x"04600001",
x"8FE40254",
x"C0001037",
x"20030020",
x"04600001",
x"200400FF",
x"C0001037",
x"2003000A",
x"04600001",
x"20060078",
x"20030003",
x"AFE20944",
x"43E2090C",
x"46000006",
x"C0000048",
x"20670000",
x"8FE20944",
x"8FE3001C",
x"43E4090C",
x"C000003F",
x"20640000",
x"AFE40910",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"20640000",
x"20C30000",
x"C000003F",
x"AFE302BC",
x"8FE602BC",
x"20030003",
x"AFE20944",
x"43E2091C",
x"46000006",
x"C0000048",
x"20670000",
x"8FE20944",
x"8FE3001C",
x"43E4091C",
x"C000003F",
x"20640000",
x"AFE40920",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE28",
x"20030003",
x"AFE20944",
x"43E2092C",
x"46000006",
x"C0000048",
x"20670000",
x"8FE20944",
x"8FE3001C",
x"43E4092C",
x"C000003F",
x"20640000",
x"AFE40930",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE2C",
x"20030003",
x"AFE20944",
x"43E2093C",
x"46000006",
x"C0000048",
x"20670000",
x"8FE20944",
x"8FE3001C",
x"43E4093C",
x"C000003F",
x"20640000",
x"AFE40940",
x"20430000",
x"20420008",
x"AC64FFFC",
x"AC670000",
x"ACC3FE30",
x"20070073",
x"C0003C7B",
x"20080003",
x"C0003CD4",
x"20030009",
x"20080000",
x"200C0000",
x"C0000081",
x"20210014",
x"200300AC",
x"C4640000",
x"44040002",
x"200300A8",
x"C4630000",
x"44030001",
x"20030004",
x"E4200010",
x"40210018",
x"C0000081",
x"20210018",
x"44000806",
x"44240802",
x"44231001",
x"20040000",
x"C4200010",
x"E4230014",
x"E4240018",
x"E421001C",
x"21830000",
x"21050000",
x"46000806",
x"46002806",
x"40210024",
x"C00039A1",
x"20210024",
x"200300A4",
x"C4650000",
x"C421001C",
x"44251000",
x"20040000",
x"20030002",
x"C4200010",
x"E4250020",
x"21050000",
x"46000806",
x"46002806",
x"40210028",
x"C00039A1",
x"20210028",
x"20030003",
x"20050001",
x"AC250024",
x"4021002C",
x"C0000081",
x"2021002C",
x"44000806",
x"C4240018",
x"44240802",
x"C4230014",
x"44231001",
x"20040000",
x"C4200010",
x"8C250024",
x"E4210028",
x"21830000",
x"46000806",
x"46002806",
x"40210030",
x"C00039A1",
x"20210030",
x"C4250020",
x"C4210028",
x"44251000",
x"20040000",
x"20080002",
x"C4200010",
x"8C250024",
x"21030000",
x"46000806",
x"46002806",
x"40210030",
x"C00039A1",
x"20210030",
x"20030002",
x"20050002",
x"AC25002C",
x"40210034",
x"C0000081",
x"20210034",
x"44000806",
x"C4240018",
x"44240802",
x"C4230014",
x"44231001",
x"20040000",
x"C4200010",
x"8C25002C",
x"E4210030",
x"21830000",
x"46000806",
x"46002806",
x"40210038",
x"C00039A1",
x"20210038",
x"C4250020",
x"C4210030",
x"44251000",
x"20040000",
x"C4200010",
x"8C25002C",
x"21030000",
x"46000806",
x"46002806",
x"40210038",
x"C00039A1",
x"20210038",
x"200A0001",
x"20090003",
x"C4200010",
x"21880000",
x"40210038",
x"C0003A9D",
x"200D0008",
x"200C0002",
x"20080004",
x"C0003B48",
x"8FEB02BC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"200C0070",
x"C0003D97",
x"20210038",
x"200D0003",
x"AC320034",
x"AC310038",
x"40210040",
x"C0003DF8",
x"C7E00134",
x"E7E002DC",
x"C7E00130",
x"E7E002D8",
x"C7E0012C",
x"E7E002D4",
x"8FE3001C",
x"40650001",
x"43E702DC",
x"43E603CC",
x"C0001D15",
x"20210040",
x"8FE3001C",
x"40660001",
x"68C000D6",
x"A0C30002",
x"03E31820",
x"8C630110",
x"8C64FFF8",
x"20050002",
x"488500CF",
x"8C64FFE4",
x"C4800000",
x"E8110002",
x"08000D8C",
x"8C65FFFC",
x"48BC0084",
x"A0CB0002",
x"8FEC06B8",
x"C4800000",
x"46206001",
x"C7E10134",
x"44205807",
x"C7EA0130",
x"45405007",
x"C7E9012C",
x"45204807",
x"216E0001",
x"20030003",
x"46000006",
x"40210040",
x"C0000048",
x"20210040",
x"20640000",
x"8FE3001C",
x"AC24003C",
x"40210044",
x"C000003F",
x"20210044",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C24003C",
x"ACA40000",
x"E4810000",
x"E48AFFFC",
x"E489FFF8",
x"8FE6001C",
x"40CD0001",
x"AC250040",
x"21A50000",
x"20660000",
x"20870000",
x"40210048",
x"C0001D15",
x"20210048",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C250040",
x"AC65FFFC",
x"AC6E0000",
x"A1840002",
x"03E42020",
x"AC8306B4",
x"218F0001",
x"216E0002",
x"C7E10130",
x"20030003",
x"46000006",
x"40210048",
x"C0000048",
x"20210048",
x"20640000",
x"8FE3001C",
x"AC240044",
x"4021004C",
x"C000003F",
x"2021004C",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240044",
x"ACA40000",
x"E48B0000",
x"E481FFFC",
x"E489FFF8",
x"8FE6001C",
x"40CD0001",
x"AC250048",
x"21A50000",
x"20660000",
x"20870000",
x"40210050",
x"C0001D15",
x"20210050",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C250048",
x"AC65FFFC",
x"AC6E0000",
x"A1E40002",
x"03E42020",
x"AC8306B4",
x"218E0002",
x"216D0003",
x"C7E1012C",
x"20030003",
x"46000006",
x"40210050",
x"C0000048",
x"20210050",
x"20640000",
x"8FE3001C",
x"AC24004C",
x"40210054",
x"C000003F",
x"20210054",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C24004C",
x"ACA40000",
x"E48B0000",
x"E48AFFFC",
x"E481FFF8",
x"8FE6001C",
x"40CB0001",
x"AC250050",
x"21650000",
x"20660000",
x"20870000",
x"40210058",
x"C0001D15",
x"20210058",
x"20430000",
x"2042000C",
x"E46CFFF8",
x"8C250050",
x"AC65FFFC",
x"AC6D0000",
x"A1C40002",
x"03E42020",
x"AC8306B4",
x"21830003",
x"AFE306B8",
x"08000D8C",
x"20040002",
x"48A40043",
x"A0C40002",
x"208C0001",
x"8FED06B8",
x"46204801",
x"8C63FFF0",
x"C7E70134",
x"C4650000",
x"44E51002",
x"C7E10130",
x"C466FFFC",
x"44260002",
x"44402000",
x"C7E2012C",
x"C460FFF8",
x"44401802",
x"44831800",
x"C42A0004",
x"45452002",
x"44832002",
x"44872801",
x"45462002",
x"44832002",
x"44812001",
x"45400002",
x"44030002",
x"44020801",
x"20030003",
x"46000006",
x"40210058",
x"C0000048",
x"20210058",
x"20640000",
x"8FE3001C",
x"AC240054",
x"4021005C",
x"C000003F",
x"2021005C",
x"20450000",
x"20420008",
x"ACA3FFFC",
x"8C240054",
x"ACA40000",
x"E4850000",
x"E484FFFC",
x"E481FFF8",
x"8FE6001C",
x"40CB0001",
x"AC250058",
x"21650000",
x"20660000",
x"20870000",
x"40210060",
x"C0001D15",
x"20210060",
x"20430000",
x"2042000C",
x"E469FFF8",
x"8C250058",
x"AC65FFFC",
x"AC6C0000",
x"A1A40002",
x"03E42020",
x"AC8306B4",
x"21A30001",
x"AFE306B8",
x"08000D8C",
x"08000D8D",
x"08000D8E",
x"20080000",
x"C7E30264",
x"8FE3025C",
x"00031822",
x"40210060",
x"C0000081",
x"20210060",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"8C300000",
x"22070000",
x"40210060",
x"C00037C4",
x"20210060",
x"200F0000",
x"20080002",
x"8FE30254",
x"69E30002",
x"08000DE2",
x"40630001",
x"AC2F005C",
x"69E30002",
x"08000DCD",
x"20040001",
x"C7E30264",
x"8FE3025C",
x"00831822",
x"40210064",
x"C0000081",
x"20210064",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"8C310038",
x"22270000",
x"40210064",
x"C00037C4",
x"20210064",
x"200E0000",
x"8C2F005C",
x"8C320034",
x"8C300000",
x"8C310038",
x"225B0000",
x"22320000",
x"23710000",
x"40210064",
x"C000383B",
x"20210064",
x"200F0001",
x"20080004",
x"8C300000",
x"8C310038",
x"8C320034",
x"22070000",
x"22500000",
x"40210064",
x"C00038AE",
x"20210064",
x"20000000",
x"0000003F",
x"EBA10037",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1001B",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA1001B",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA1000D",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"443D0801",
x"EBA10006",
x"E8300003",
x"44200006",
x"E0000000",
x"443D0800",
x"08000DE4",
x"443D0801",
x"08000DE4",
x"04002000",
x"20030030",
x"68830007",
x"20030039",
x"68640003",
x"20030000",
x"08000E56",
x"20030001",
x"08000E58",
x"20030001",
x"48600037",
x"8FE30008",
x"48600009",
x"2003002D",
x"48A30004",
x"2003FFFF",
x"AFE30008",
x"08000E62",
x"20030001",
x"AFE30008",
x"08000E63",
x"8FE30004",
x"A0650003",
x"A0630001",
x"00A32820",
x"40830030",
x"00A31820",
x"AFE30004",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000E72",
x"20030001",
x"08000E74",
x"20030001",
x"48600014",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08000E7E",
x"20030001",
x"AFE30008",
x"08000E7F",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"08000E4E",
x"8FE30008",
x"487C0003",
x"8FE30004",
x"E0000000",
x"8FE30004",
x"00031822",
x"E0000000",
x"48C00021",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000E98",
x"20030001",
x"08000E9A",
x"20030001",
x"48600014",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08000EA4",
x"20030001",
x"AFE30008",
x"08000EA5",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"08000E4E",
x"20060000",
x"08000E4E",
x"8FE30008",
x"487C0003",
x"8FE30004",
x"E0000000",
x"8FE30004",
x"00031822",
x"E0000000",
x"04002000",
x"20030030",
x"68830007",
x"20030039",
x"68640003",
x"20030000",
x"08000EBF",
x"20030001",
x"08000EC1",
x"20030001",
x"48600032",
x"8FE30018",
x"48600009",
x"2003002D",
x"48A30004",
x"2003FFFF",
x"AFE30018",
x"08000ECB",
x"20030001",
x"AFE30018",
x"08000ECC",
x"8FE3000C",
x"A0650003",
x"A0630001",
x"00A32820",
x"40830030",
x"00A31820",
x"AFE3000C",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000EDB",
x"20030001",
x"08000EDD",
x"20030001",
x"48600014",
x"8FE30018",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30018",
x"08000EE7",
x"20030001",
x"AFE30018",
x"08000EE8",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"08000EB7",
x"20A30000",
x"E0000000",
x"48C00021",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08000EFC",
x"20030001",
x"08000EFE",
x"20030001",
x"48600014",
x"8FE30018",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30018",
x"08000F08",
x"20030001",
x"AFE30018",
x"08000F09",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"08000EB7",
x"20060000",
x"08000EB7",
x"20830000",
x"E0000000",
x"04001800",
x"20050030",
x"68650007",
x"20050039",
x"68A30003",
x"20050000",
x"08000F1E",
x"20050001",
x"08000F20",
x"20050001",
x"48A00027",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000F35",
x"20040001",
x"08000F37",
x"20040001",
x"4880000F",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"08000F16",
x"E0000000",
x"4880001C",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08000F50",
x"20040001",
x"08000F52",
x"20040001",
x"4880000F",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"08000F16",
x"20040000",
x"08000F16",
x"E0000000",
x"012A1820",
x"A8650001",
x"00A63818",
x"01491822",
x"6B830003",
x"21230000",
x"E0000000",
x"68E40068",
x"48E40003",
x"20A30000",
x"E0000000",
x"01251820",
x"A8670001",
x"00E64018",
x"00A91822",
x"6B830003",
x"21230000",
x"E0000000",
x"69040030",
x"49040003",
x"20E30000",
x"E0000000",
x"01271820",
x"A8680001",
x"01062818",
x"00E91822",
x"6B830003",
x"21230000",
x"E0000000",
x"68A40014",
x"48A40003",
x"21030000",
x"E0000000",
x"01281820",
x"A8650001",
x"00A63818",
x"01091822",
x"6B830003",
x"21230000",
x"E0000000",
x"68E40006",
x"48E40003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"08000F64",
x"210A0000",
x"20A90000",
x"08000F64",
x"01071820",
x"A8650001",
x"00A64818",
x"00E81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"21090000",
x"08000F64",
x"20EA0000",
x"20A90000",
x"08000F64",
x"00E51820",
x"A8680001",
x"01064818",
x"00A71822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240015",
x"49240003",
x"21030000",
x"E0000000",
x"00E81820",
x"A8650001",
x"00A64818",
x"01071822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000F64",
x"210A0000",
x"20A90000",
x"08000F64",
x"01051820",
x"A8670001",
x"00E64818",
x"00A81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20E30000",
x"E0000000",
x"20EA0000",
x"21090000",
x"08000F64",
x"20AA0000",
x"20E90000",
x"08000F64",
x"00AA1820",
x"A8680001",
x"01063818",
x"01451822",
x"6B830003",
x"20A30000",
x"E0000000",
x"68E40031",
x"48E40003",
x"21030000",
x"E0000000",
x"00A81820",
x"A8670001",
x"00E64818",
x"01051822",
x"6B830003",
x"20A30000",
x"E0000000",
x"69240015",
x"49240003",
x"20E30000",
x"E0000000",
x"00A71820",
x"A8680001",
x"01064818",
x"00E51822",
x"6B830003",
x"20A30000",
x"E0000000",
x"69240007",
x"49240003",
x"21030000",
x"E0000000",
x"210A0000",
x"20A90000",
x"08000F64",
x"20EA0000",
x"21090000",
x"08000F64",
x"00E81820",
x"A8650001",
x"00A64818",
x"01071822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000F64",
x"210A0000",
x"20A90000",
x"08000F64",
x"010A1820",
x"A8670001",
x"00E62818",
x"01481822",
x"6B830003",
x"21030000",
x"E0000000",
x"68A40015",
x"48A40003",
x"20E30000",
x"E0000000",
x"01071820",
x"A8650001",
x"00A64818",
x"00E81822",
x"6B830003",
x"21030000",
x"E0000000",
x"69240007",
x"49240003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"21090000",
x"08000F64",
x"20EA0000",
x"20A90000",
x"08000F64",
x"00EA1820",
x"A8650001",
x"00A64018",
x"01471822",
x"6B830003",
x"20E30000",
x"E0000000",
x"69040007",
x"49040003",
x"20A30000",
x"E0000000",
x"20AA0000",
x"20E90000",
x"08000F64",
x"20A90000",
x"08000F64",
x"200303E8",
x"68830002",
x"E0000000",
x"688000CF",
x"20060064",
x"200C0000",
x"200A000A",
x"20090005",
x"200501F4",
x"AC240000",
x"68A4002D",
x"48A40003",
x"20030005",
x"0800106D",
x"200B0002",
x"200500C8",
x"68A40015",
x"48A40003",
x"20030002",
x"0800105B",
x"20090001",
x"20050064",
x"68A4000A",
x"48A40003",
x"20030001",
x"08001056",
x"212A0000",
x"21890000",
x"40210008",
x"C0000F64",
x"20210008",
x"0800105B",
x"216A0000",
x"40210008",
x"C0000F64",
x"20210008",
x"0800106D",
x"200A0003",
x"2005012C",
x"68A40009",
x"48A40003",
x"20030003",
x"08001066",
x"21690000",
x"40210008",
x"C0000F64",
x"20210008",
x"0800106D",
x"215B0000",
x"212A0000",
x"23690000",
x"40210008",
x"C0000F64",
x"20210008",
x"08001093",
x"200B0007",
x"200502BC",
x"68A40014",
x"48A40003",
x"20030007",
x"08001083",
x"200A0006",
x"20050258",
x"68A40008",
x"48A40003",
x"20030006",
x"0800107D",
x"40210008",
x"C0000F64",
x"20210008",
x"08001083",
x"21490000",
x"216A0000",
x"40210008",
x"C0000F64",
x"20210008",
x"08001093",
x"20090008",
x"20050320",
x"68A4000A",
x"48A40003",
x"20030008",
x"0800108F",
x"212A0000",
x"21690000",
x"40210008",
x"C0000F64",
x"20210008",
x"08001093",
x"40210008",
x"C0000F64",
x"20210008",
x"60650064",
x"8C240000",
x"00852022",
x"68030003",
x"200D0000",
x"0800109D",
x"20050030",
x"00A31820",
x"04600001",
x"200D0001",
x"2006000A",
x"200C0000",
x"200A000A",
x"20090005",
x"20050032",
x"AC240004",
x"68A4002D",
x"48A40003",
x"20030005",
x"080010CF",
x"200B0002",
x"20050014",
x"68A40015",
x"48A40003",
x"20030002",
x"080010BD",
x"20090001",
x"2005000A",
x"68A4000A",
x"48A40003",
x"20030001",
x"080010B8",
x"212A0000",
x"21890000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010BD",
x"216A0000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010CF",
x"200A0003",
x"2005001E",
x"68A40009",
x"48A40003",
x"20030003",
x"080010C8",
x"21690000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010CF",
x"215B0000",
x"212A0000",
x"23690000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010F5",
x"200B0007",
x"20050046",
x"68A40014",
x"48A40003",
x"20030007",
x"080010E5",
x"200A0006",
x"2005003C",
x"68A40008",
x"48A40003",
x"20030006",
x"080010DF",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010E5",
x"21490000",
x"216A0000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010F5",
x"20090008",
x"20050050",
x"68A4000A",
x"48A40003",
x"20030008",
x"080010F1",
x"212A0000",
x"21690000",
x"4021000C",
x"C0000F64",
x"2021000C",
x"080010F5",
x"4021000C",
x"C0000F64",
x"2021000C",
x"6065000A",
x"8C240004",
x"00852022",
x"68030009",
x"49A00003",
x"20050000",
x"08001100",
x"20050030",
x"00A31820",
x"04600001",
x"20050001",
x"08001105",
x"20050030",
x"00A31820",
x"04600001",
x"20050001",
x"20030030",
x"00641820",
x"04600001",
x"E0000000",
x"2003002D",
x"04600001",
x"00042022",
x"08001037",
x"2003003C",
x"6A030002",
x"E0000000",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200E0030",
x"68AE0007",
x"200E0039",
x"69C50003",
x"200E0000",
x"0800111C",
x"200E0001",
x"0800111E",
x"200E0001",
x"49C00013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001124",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206E0000",
x"08001136",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206E0000",
x"49DD0003",
x"20030000",
x"08001AF2",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200B0030",
x"68AB0007",
x"200B0039",
x"69650003",
x"200B0000",
x"08001145",
x"200B0001",
x"08001147",
x"200B0001",
x"49600013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"0800114D",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206B0000",
x"0800115F",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206B0000",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200F0030",
x"68AF0007",
x"200F0039",
x"69E50003",
x"200F0000",
x"0800116B",
x"200F0001",
x"0800116D",
x"200F0001",
x"49E00013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001173",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206F0000",
x"08001185",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206F0000",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200D0030",
x"68AD0007",
x"200D0039",
x"69A50003",
x"200D0000",
x"08001191",
x"200D0001",
x"08001193",
x"200D0001",
x"49A00013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001199",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206D0000",
x"080011AB",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206D0000",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20680000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080011C1",
x"20030001",
x"080011C3",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080011C9",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080011D9",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080011E3",
x"20040001",
x"080011E5",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080011FB",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"0800120C",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08001211",
x"44000807",
x"E5010000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08001222",
x"20030001",
x"08001224",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"0800122A",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"0800123A",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08001244",
x"20040001",
x"08001246",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"0800125C",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"0800126D",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08001272",
x"44000807",
x"E501FFFC",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08001283",
x"20030001",
x"08001285",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"0800128B",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"0800129B",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080012A5",
x"20040001",
x"080012A7",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080012BD",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"080012CE",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080012D3",
x"44000807",
x"E501FFF8",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"206C0000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080012EA",
x"20030001",
x"080012EC",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080012F2",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001302",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800130C",
x"20040001",
x"0800130E",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001324",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08001335",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800133A",
x"44000807",
x"E5810000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800134B",
x"20030001",
x"0800134D",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08001353",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001363",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800136D",
x"20040001",
x"0800136F",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001385",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08001396",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800139B",
x"44000807",
x"E581FFFC",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080013AC",
x"20030001",
x"080013AE",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080013B4",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080013C4",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080013CE",
x"20040001",
x"080013D0",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080013E6",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"080013F7",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080013FC",
x"44000807",
x"E581FFF8",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800140D",
x"20030001",
x"0800140F",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08001415",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001425",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800142F",
x"20040001",
x"08001431",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001447",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002006",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44800000",
x"08001458",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44002006",
x"0800145D",
x"44002007",
x"20030002",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"206A0000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08001473",
x"20030001",
x"08001475",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"0800147B",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"0800148B",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08001495",
x"20040001",
x"08001497",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080014AD",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"080014BE",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080014C3",
x"44000807",
x"E5410000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080014D4",
x"20030001",
x"080014D6",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080014DC",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080014EC",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080014F6",
x"20040001",
x"080014F8",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"0800150E",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"0800151F",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"08001524",
x"44000807",
x"E541FFFC",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20690000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800153B",
x"20030001",
x"0800153D",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08001543",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001553",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800155D",
x"20040001",
x"0800155F",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001575",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"08001586",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800158B",
x"44000807",
x"E5210000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800159C",
x"20030001",
x"0800159E",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080015A4",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080015B4",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080015BE",
x"20040001",
x"080015C0",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080015D6",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"080015E7",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080015EC",
x"44000807",
x"E521FFFC",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080015FD",
x"20030001",
x"080015FF",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08001605",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001615",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800161F",
x"20040001",
x"08001621",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001637",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"08001648",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800164D",
x"44000807",
x"E521FFF8",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20670000",
x"49A00002",
x"0800177E",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08001666",
x"20030001",
x"08001668",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"0800166E",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"0800167E",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"08001688",
x"20040001",
x"0800168A",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"080016A0",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44002806",
x"8FE30010",
x"C0000081",
x"44001806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44600003",
x"44A00000",
x"080016B1",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"080016B6",
x"44000807",
x"200300CC",
x"C4630000",
x"44230002",
x"E4E00000",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"080016CA",
x"20030001",
x"080016CC",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"080016D2",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"080016E2",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"080016EC",
x"20040001",
x"080016EE",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001704",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44003006",
x"8FE30010",
x"C0000081",
x"44002806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44A00003",
x"44C00000",
x"08001715",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800171A",
x"44000807",
x"44230002",
x"E4E0FFFC",
x"20030000",
x"AFE3000C",
x"20030000",
x"AFE30010",
x"20030001",
x"AFE30014",
x"20030000",
x"AFE30018",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"0800172C",
x"20030001",
x"0800172E",
x"20030001",
x"48600012",
x"8FE30018",
x"48600004",
x"20030001",
x"AFE30018",
x"08001734",
x"8FE3000C",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE3000C",
x"20060001",
x"40210004",
x"C0000EB7",
x"20210004",
x"08001744",
x"20060000",
x"40210004",
x"C0000EB7",
x"20210004",
x"2004002E",
x"4864002E",
x"04001800",
x"20040030",
x"68640007",
x"20040039",
x"68830003",
x"20040000",
x"0800174E",
x"20040001",
x"08001750",
x"20040001",
x"48800012",
x"8FE40010",
x"A0850003",
x"A0840001",
x"00A42020",
x"40630030",
x"00831820",
x"AFE30010",
x"8FE30014",
x"A0640003",
x"A0630001",
x"00831820",
x"AFE30014",
x"20040001",
x"40210004",
x"C0000F16",
x"20210004",
x"08001766",
x"20040000",
x"40210004",
x"C0000F16",
x"20210004",
x"8FE3000C",
x"40210004",
x"C0000081",
x"44003006",
x"8FE30010",
x"C0000081",
x"44002806",
x"8FE30014",
x"C0000081",
x"20210004",
x"44A00003",
x"44C00000",
x"08001777",
x"8FE3000C",
x"40210004",
x"C0000081",
x"20210004",
x"8FE30018",
x"487C0003",
x"44000806",
x"0800177C",
x"44000807",
x"44230002",
x"E4E0FFF8",
x"20050002",
x"49650003",
x"20050001",
x"08001786",
x"E8900003",
x"20050000",
x"08001786",
x"20050001",
x"20030004",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20640000",
x"20430000",
x"2042002C",
x"AC64FFD8",
x"AC67FFDC",
x"AC69FFE0",
x"AC6AFFE4",
x"AC65FFE8",
x"AC6CFFEC",
x"AC68FFF0",
x"AC6DFFF4",
x"AC6FFFF8",
x"AC6BFFFC",
x"AC6E0000",
x"A2040002",
x"03E42020",
x"AC830110",
x"20030003",
x"49630032",
x"C5010000",
x"C830000D",
x"C8300008",
x"EA010004",
x"200300A0",
x"C4600000",
x"080017A7",
x"200300C8",
x"C4600000",
x"080017A9",
x"46000006",
x"44210802",
x"44010003",
x"080017AD",
x"46000006",
x"E5000000",
x"C501FFFC",
x"C830000D",
x"C8300008",
x"EA010004",
x"200300A0",
x"C4600000",
x"080017B7",
x"200300C8",
x"C4600000",
x"080017B9",
x"46000006",
x"44210802",
x"44010003",
x"080017BD",
x"46000006",
x"E500FFFC",
x"C501FFF8",
x"C830000D",
x"C8300008",
x"EA010004",
x"200300A0",
x"C4600000",
x"080017C7",
x"200300C8",
x"C4600000",
x"080017C9",
x"46000006",
x"44210802",
x"44010003",
x"080017CD",
x"46000006",
x"E500FFF8",
x"080017EB",
x"20030002",
x"4963001B",
x"C5010000",
x"44211002",
x"C500FFFC",
x"44000002",
x"44401000",
x"C500FFF8",
x"44000002",
x"44400000",
x"44001004",
x"C8500006",
x"E8900003",
x"46820003",
x"080017DF",
x"46220003",
x"080017E2",
x"200300C8",
x"C4600000",
x"44200802",
x"E5010000",
x"C501FFFC",
x"44200802",
x"E501FFFC",
x"C501FFF8",
x"44200002",
x"E500FFF8",
x"080017EB",
x"49A00002",
x"08001AF1",
x"C4E30000",
x"46C31001",
x"200300F0",
x"C4640000",
x"200300EC",
x"C46E0000",
x"E8500003",
x"44400806",
x"080017F7",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"0800181D",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800180E",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001809",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"0800180E",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"0800181D",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001818",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"0800181D",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08001840",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001831",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800182C",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08001831",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08001840",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800183B",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08001840",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8800006",
x"EA020003",
x"20030000",
x"08001845",
x"20030001",
x"0800184A",
x"EA020003",
x"20030001",
x"0800184A",
x"20030000",
x"E8800003",
x"44000806",
x"0800184E",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001852",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44007807",
x"08001865",
x"44007806",
x"E8700003",
x"44600806",
x"08001869",
x"44600807",
x"E42F0000",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001890",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001881",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800187C",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001881",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001890",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800188B",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001890",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"080018B3",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080018A4",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"0800189F",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080018A4",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"080018B3",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080018AE",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080018B3",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8800006",
x"EA030003",
x"20030000",
x"080018B8",
x"20030001",
x"080018BD",
x"EA030003",
x"20030001",
x"080018BD",
x"20030000",
x"E8800003",
x"44000806",
x"080018C1",
x"47A00801",
x"EAC10003",
x"44200006",
x"080018C5",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44003807",
x"080018D8",
x"44003806",
x"C4E3FFFC",
x"46C31001",
x"E8500003",
x"44400806",
x"080018DE",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001904",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080018F5",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080018F0",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080018F5",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001904",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080018FF",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001904",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001927",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001918",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001913",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001918",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001927",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001922",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001927",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8800006",
x"EA020003",
x"20030000",
x"0800192C",
x"20030001",
x"08001931",
x"EA020003",
x"20030001",
x"08001931",
x"20030000",
x"E8800003",
x"44000806",
x"08001935",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001939",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200803",
x"45C10002",
x"44210802",
x"46210800",
x"44010003",
x"48600003",
x"44006807",
x"0800194C",
x"44006806",
x"E8700003",
x"44600806",
x"08001950",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001976",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001967",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001962",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001967",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001976",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001971",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001976",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001999",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800198A",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001985",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"0800198A",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001999",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001994",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001999",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8800006",
x"EA030003",
x"20030000",
x"0800199E",
x"20030001",
x"080019A3",
x"EA030003",
x"20030001",
x"080019A3",
x"20030000",
x"E8800003",
x"44000806",
x"080019A7",
x"47A00801",
x"EAC10003",
x"44200006",
x"080019AB",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200803",
x"45C10002",
x"44210802",
x"46210800",
x"44010003",
x"48600003",
x"44004807",
x"080019BE",
x"44004806",
x"C4E3FFF8",
x"46C31001",
x"E8500003",
x"44400806",
x"080019C4",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"080019EA",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"080019DB",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080019D6",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080019DB",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"080019EA",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"080019E5",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080019EA",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A0D",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"080019FE",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"080019F9",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"080019FE",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A0D",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001A08",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A0D",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8800006",
x"EA020003",
x"20030000",
x"08001A12",
x"20030001",
x"08001A17",
x"EA020003",
x"20030001",
x"08001A17",
x"20030000",
x"E8800003",
x"44000806",
x"08001A1B",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001A1F",
x"44810001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44001007",
x"08001A32",
x"44001006",
x"E8700003",
x"44600806",
x"08001A36",
x"44600807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08001A5C",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001A4D",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001A48",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A4D",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A5C",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001A57",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A5C",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A7F",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08001A70",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001A6B",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A70",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A7F",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08001A7A",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08001A7F",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8800006",
x"EA030003",
x"20030000",
x"08001A84",
x"20030001",
x"08001A89",
x"EA030003",
x"20030001",
x"08001A89",
x"20030000",
x"E8800003",
x"44000806",
x"08001A8D",
x"47A00801",
x"EAC10003",
x"44200006",
x"08001A91",
x"44810001",
x"44150802",
x"44210002",
x"44191803",
x"47431801",
x"44031803",
x"47031801",
x"44031803",
x"46E31801",
x"44030003",
x"46200001",
x"44200003",
x"45C00802",
x"44000002",
x"46200000",
x"44200803",
x"48600003",
x"44200007",
x"08001AA4",
x"44200006",
x"45A26002",
x"44E92802",
x"44A21802",
x"C42F0000",
x"45E00802",
x"44615001",
x"45E90802",
x"44222002",
x"44E01802",
x"44833000",
x"45A05802",
x"44A02002",
x"45E21802",
x"44834000",
x"44200802",
x"44E20002",
x"44202801",
x"45204807",
x"44ED3802",
x"45ED2002",
x"C5000000",
x"C502FFFC",
x"C503FFF8",
x"458C0802",
x"44016802",
x"456B0802",
x"44410802",
x"45A16800",
x"45290802",
x"44610802",
x"45A10800",
x"E5010000",
x"454A0802",
x"44016802",
x"45080802",
x"44410802",
x"45A16800",
x"44E70802",
x"44610802",
x"45A10800",
x"E501FFFC",
x"44C60802",
x"44016802",
x"44A50802",
x"44410802",
x"45A16800",
x"44840802",
x"44610802",
x"45A10800",
x"E501FFF8",
x"440A0802",
x"44266802",
x"44480802",
x"44250802",
x"45A16800",
x"44670802",
x"44240802",
x"45A10800",
x"45C10802",
x"E4E10000",
x"440C0802",
x"44263002",
x"444B0002",
x"44051002",
x"44C22800",
x"44691802",
x"44641002",
x"44A21000",
x"45C21002",
x"E4E2FFFC",
x"442A0802",
x"44080002",
x"44200800",
x"44670002",
x"44200000",
x"45C00002",
x"E4E0FFF8",
x"20030001",
x"48600003",
x"AFF0001C",
x"E0000000",
x"22100001",
x"0800110D",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002000",
x"20070030",
x"68870007",
x"20070039",
x"68E40003",
x"20070000",
x"08001B03",
x"20070001",
x"08001B05",
x"20070001",
x"48E00036",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001B0B",
x"8FE30004",
x"A0650003",
x"A0630001",
x"00A32820",
x"40830030",
x"00A31820",
x"AFE30004",
x"04002800",
x"20070030",
x"68A70007",
x"20070039",
x"68E50003",
x"20070000",
x"08001B1A",
x"20070001",
x"08001B1C",
x"20070001",
x"48E00018",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08001B26",
x"20030001",
x"AFE30008",
x"08001B27",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"20670000",
x"08001B3A",
x"8FE70008",
x"48FC0003",
x"8FE70004",
x"08001B3A",
x"8FE70004",
x"00073822",
x"08001B62",
x"04002800",
x"20070030",
x"68A70007",
x"20070039",
x"68E50003",
x"20070000",
x"08001B43",
x"20070001",
x"08001B45",
x"20070001",
x"48E00018",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08001B4F",
x"20030001",
x"AFE30008",
x"08001B50",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"20670000",
x"08001B62",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"20670000",
x"48FD0004",
x"21030001",
x"2004FFFF",
x"0800003F",
x"21090001",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"20040030",
x"68A40007",
x"20040039",
x"68850003",
x"20040000",
x"08001B73",
x"20040001",
x"08001B75",
x"20040001",
x"48800013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001B7B",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"20640000",
x"08001B8D",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"20640000",
x"AC270000",
x"AC280004",
x"489D0007",
x"21230001",
x"2004FFFF",
x"4021000C",
x"C000003F",
x"2021000C",
x"08001BA1",
x"21230001",
x"AC240008",
x"AC29000C",
x"20680000",
x"40210014",
x"C0001AF7",
x"20210014",
x"8C29000C",
x"A1250002",
x"8C240008",
x"6C652000",
x"8C280004",
x"A1040002",
x"8C270000",
x"6C643800",
x"E0000000",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"20030030",
x"68A30007",
x"20030039",
x"68650003",
x"20030000",
x"08001BB2",
x"20030001",
x"08001BB4",
x"20030001",
x"48600012",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001BBA",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"08001BCA",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"487D0008",
x"20030001",
x"2004FFFF",
x"40210004",
x"C000003F",
x"20210004",
x"20650000",
x"08001BDA",
x"20080001",
x"AC230000",
x"40210008",
x"C0001AF7",
x"20210008",
x"20650000",
x"8C230000",
x"ACA30000",
x"8CA30000",
x"487D0004",
x"21630001",
x"20A40000",
x"0800003F",
x"216A0001",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04003800",
x"20030030",
x"68E30007",
x"20030039",
x"68670003",
x"20030000",
x"08001BEC",
x"20030001",
x"08001BEE",
x"20030001",
x"AC250004",
x"48600013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001BF5",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40E30030",
x"00831820",
x"AFE30004",
x"20060001",
x"20E50000",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"08001C07",
x"20060000",
x"20E50000",
x"4021000C",
x"C0000E4E",
x"2021000C",
x"487D0008",
x"20030001",
x"2004FFFF",
x"4021000C",
x"C000003F",
x"2021000C",
x"20640000",
x"08001C17",
x"20080001",
x"AC230008",
x"40210010",
x"C0001AF7",
x"20210010",
x"20640000",
x"8C230008",
x"AC830000",
x"8C830000",
x"AC2B000C",
x"487D0006",
x"21430001",
x"40210014",
x"C000003F",
x"20210014",
x"08001C2A",
x"21430001",
x"AC240010",
x"AC2A0014",
x"206B0000",
x"4021001C",
x"C0001BA6",
x"2021001C",
x"8C2A0014",
x"A1460002",
x"8C240010",
x"6C662000",
x"8C2B000C",
x"A1640002",
x"8C250004",
x"6C642800",
x"E0000000",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002000",
x"200A0030",
x"688A0007",
x"200A0039",
x"69440003",
x"200A0000",
x"08001C3B",
x"200A0001",
x"08001C3D",
x"200A0001",
x"49400036",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001C43",
x"8FE30004",
x"A0650003",
x"A0630001",
x"00A32820",
x"40830030",
x"00A31820",
x"AFE30004",
x"04002800",
x"200A0030",
x"68AA0007",
x"200A0039",
x"69450003",
x"200A0000",
x"08001C52",
x"200A0001",
x"08001C54",
x"200A0001",
x"49400018",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08001C5E",
x"20030001",
x"AFE30008",
x"08001C5F",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206A0000",
x"08001C72",
x"8FEA0008",
x"495C0003",
x"8FEA0004",
x"08001C72",
x"8FEA0004",
x"000A5022",
x"08001C9A",
x"04002800",
x"200A0030",
x"68AA0007",
x"200A0039",
x"69450003",
x"200A0000",
x"08001C7B",
x"200A0001",
x"08001C7D",
x"200A0001",
x"49400018",
x"8FE30008",
x"48600009",
x"2003002D",
x"48830004",
x"2003FFFF",
x"AFE30008",
x"08001C87",
x"20030001",
x"AFE30008",
x"08001C88",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206A0000",
x"08001C9A",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206A0000",
x"495D0007",
x"20030001",
x"2004FFFF",
x"40210004",
x"C000003F",
x"20210004",
x"08001CD4",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200C0030",
x"68AC0007",
x"200C0039",
x"69850003",
x"200C0000",
x"08001CAD",
x"200C0001",
x"08001CAF",
x"200C0001",
x"49800013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001CB5",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206C0000",
x"08001CC7",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206C0000",
x"499D0007",
x"20030002",
x"2004FFFF",
x"40210004",
x"C000003F",
x"20210004",
x"08001CD3",
x"20080002",
x"40210004",
x"C0001AF7",
x"20210004",
x"AC6CFFFC",
x"AC6A0000",
x"8C640000",
x"489D0002",
x"E0000000",
x"A1640002",
x"03E42020",
x"AC830200",
x"216B0001",
x"20030000",
x"AFE30004",
x"20030000",
x"AFE30008",
x"04002800",
x"200A0030",
x"68AA0007",
x"200A0039",
x"69450003",
x"200A0000",
x"08001CE7",
x"200A0001",
x"08001CE9",
x"200A0001",
x"49400013",
x"8FE30008",
x"48600004",
x"20030001",
x"AFE30008",
x"08001CEF",
x"8FE30004",
x"A0640003",
x"A0630001",
x"00832020",
x"40A30030",
x"00831820",
x"AFE30004",
x"20060001",
x"40210004",
x"C0000E4E",
x"20210004",
x"206A0000",
x"08001D01",
x"20060000",
x"40210004",
x"C0000E4E",
x"20210004",
x"206A0000",
x"495D0007",
x"20030001",
x"2004FFFF",
x"40210004",
x"C000003F",
x"20210004",
x"08001D0D",
x"20080001",
x"40210004",
x"C0001AF7",
x"20210004",
x"AC6A0000",
x"8C640000",
x"489D0002",
x"E0000000",
x"A1640002",
x"03E42020",
x"AC830200",
x"216B0001",
x"08001C2F",
x"68A000C6",
x"A0A30002",
x"03E31820",
x"8C690110",
x"8D23FFFC",
x"487C0042",
x"20030006",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E00000",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"08001D27",
x"200A0001",
x"8D28FFF0",
x"C5010000",
x"488A0003",
x"44200007",
x"08001D2D",
x"44200006",
x"E4600000",
x"C4E00000",
x"46200003",
x"E460FFFC",
x"08001D33",
x"E470FFFC",
x"C4E0FFFC",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"08001D3A",
x"200A0001",
x"8D28FFF0",
x"C501FFFC",
x"488A0003",
x"44200007",
x"08001D40",
x"44200006",
x"E460FFF8",
x"C4E0FFFC",
x"46200003",
x"E460FFF4",
x"08001D46",
x"E470FFF4",
x"C4E0FFF8",
x"C8100011",
x"8D24FFE8",
x"E8100003",
x"200A0000",
x"08001D4D",
x"200A0001",
x"8D28FFF0",
x"C501FFF8",
x"488A0003",
x"44200007",
x"08001D53",
x"44200006",
x"E460FFF0",
x"C4E0FFF8",
x"46200003",
x"E460FFEC",
x"08001D59",
x"E470FFEC",
x"A0A40002",
x"6CC41800",
x"08001DD9",
x"20040002",
x"48640026",
x"20030004",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E10000",
x"8D24FFF0",
x"C4800000",
x"44201002",
x"C4E1FFFC",
x"C480FFFC",
x"44200002",
x"44401000",
x"C4E1FFF8",
x"C480FFF8",
x"44200002",
x"44400000",
x"EA000003",
x"E4700000",
x"08001D80",
x"46800803",
x"E4610000",
x"C4810000",
x"44200803",
x"44200807",
x"E461FFFC",
x"C481FFFC",
x"44200803",
x"44200807",
x"E461FFF8",
x"C481FFF8",
x"44200003",
x"44000007",
x"E460FFF4",
x"A0A40002",
x"6CC41800",
x"08001DD9",
x"20030005",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"C4E00000",
x"C4E1FFFC",
x"C4E2FFF8",
x"44001802",
x"8D24FFF0",
x"C4850000",
x"44652002",
x"44211802",
x"C486FFFC",
x"44661802",
x"44833800",
x"44421802",
x"C484FFF8",
x"44641802",
x"44E33800",
x"8D28FFF4",
x"49000003",
x"44E01806",
x"08001DA8",
x"44224002",
x"8D24FFDC",
x"C4830000",
x"45031802",
x"44E34000",
x"44403802",
x"C483FFFC",
x"44E31802",
x"45034000",
x"44013802",
x"C483FFF8",
x"44E31802",
x"45031800",
x"44050002",
x"44000007",
x"44260802",
x"44200807",
x"44441002",
x"44401007",
x"E4630000",
x"49000005",
x"E460FFFC",
x"E461FFF8",
x"E462FFF4",
x"08001DD3",
x"C4E5FFF8",
x"8D24FFDC",
x"C484FFFC",
x"44A43002",
x"C4E5FFFC",
x"C484FFF8",
x"44A42002",
x"44C42000",
x"44952002",
x"44040001",
x"E460FFFC",
x"C4E4FFF8",
x"C4800000",
x"44802802",
x"C4E40000",
x"C480FFF8",
x"44800002",
x"44A00000",
x"44150002",
x"44200001",
x"E460FFF8",
x"C4E1FFFC",
x"C4800000",
x"44202002",
x"C4E10000",
x"C480FFFC",
x"44200002",
x"44800000",
x"44150002",
x"44400001",
x"E460FFF4",
x"C8700004",
x"46230003",
x"E460FFF0",
x"08001DD7",
x"A0A40002",
x"6CC41800",
x"40A50001",
x"08001D15",
x"E0000000",
x"6880009C",
x"A0850002",
x"03E52820",
x"8CA50110",
x"8CA8FFD8",
x"8CA7FFFC",
x"C4610000",
x"8CA6FFEC",
x"C4C00000",
x"44200001",
x"E5000000",
x"C461FFFC",
x"C4C0FFFC",
x"44200001",
x"E500FFFC",
x"C461FFF8",
x"C4C0FFF8",
x"44200001",
x"E500FFF8",
x"20060002",
x"48E6000F",
x"8CA5FFF0",
x"C5010000",
x"C503FFFC",
x"C502FFF8",
x"C4A00000",
x"44010802",
x"C4A0FFFC",
x"44030002",
x"44200800",
x"C4A0FFF8",
x"44020002",
x"44200000",
x"E500FFF4",
x"08001E28",
x"20060002",
x"68C70002",
x"08001E28",
x"C5020000",
x"C501FFFC",
x"C500FFF8",
x"44422002",
x"8CA6FFF0",
x"C4C30000",
x"44832802",
x"44212002",
x"C4C3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4C3FFF8",
x"44831802",
x"44A32000",
x"8CA6FFF4",
x"48C00003",
x"44801806",
x"08001E22",
x"44202802",
x"8CA5FFDC",
x"C4A30000",
x"44A31802",
x"44832000",
x"44021802",
x"C4A0FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C4A0FFF8",
x"44201802",
x"44831800",
x"20050003",
x"48E50003",
x"44710001",
x"08001E27",
x"44600006",
x"E500FFF4",
x"40880001",
x"6900004E",
x"A1040002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C4610000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C461FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C461FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08001E75",
x"20050002",
x"68A60002",
x"08001E75",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08001E6F",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08001E74",
x"44600006",
x"E4E0FFF4",
x"41040001",
x"08001DDC",
x"E0000000",
x"E0000000",
x"A0A30002",
x"4C833000",
x"48DD0003",
x"20030001",
x"E0000000",
x"A0C30002",
x"03E31820",
x"8C670110",
x"8CE3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CE6FFFC",
x"48DC0024",
x"E8100003",
x"44003006",
x"08001E8E",
x"44003007",
x"8CE3FFF0",
x"C4600000",
x"E8C00003",
x"20060000",
x"08001EA4",
x"E8500003",
x"44400006",
x"08001E97",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20060000",
x"08001EA4",
x"E8300003",
x"44200006",
x"08001E9F",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20060000",
x"08001EA4",
x"20060001",
x"48C00007",
x"8CE3FFE8",
x"48600003",
x"20030001",
x"08001EAA",
x"20030000",
x"08001EAC",
x"8CE3FFE8",
x"08001EED",
x"20030002",
x"48C30014",
x"8CE3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CE3FFE8",
x"E8100003",
x"20060000",
x"08001EBD",
x"20060001",
x"48660003",
x"20030001",
x"08001EC1",
x"20030000",
x"08001EED",
x"44003802",
x"8CE3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CE3FFF4",
x"48600003",
x"44E03006",
x"08001EDF",
x"44414002",
x"8CE3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48C30003",
x"44D10001",
x"08001EE4",
x"44C00006",
x"8CE3FFE8",
x"E8100003",
x"20060000",
x"08001EE9",
x"20060001",
x"48660003",
x"20030001",
x"08001EED",
x"20030000",
x"4860007B",
x"20A70001",
x"A0E30002",
x"4C832800",
x"48BD0003",
x"20030001",
x"E0000000",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08001F04",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"08001F1A",
x"E8500003",
x"44400006",
x"08001F0D",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"08001F1A",
x"E8300003",
x"44200006",
x"08001F15",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"08001F1A",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08001F20",
x"20030000",
x"08001F22",
x"8CC3FFE8",
x"08001F63",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001F33",
x"20050001",
x"48650003",
x"20030001",
x"08001F37",
x"20030000",
x"08001F63",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"08001F55",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"08001F5A",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08001F5F",
x"20050001",
x"48650003",
x"20030001",
x"08001F63",
x"20030000",
x"48600003",
x"20E50001",
x"08001E79",
x"20030000",
x"E0000000",
x"20030000",
x"E0000000",
x"A1030002",
x"4C834800",
x"493D0003",
x"20030000",
x"E0000000",
x"A1230002",
x"03E31820",
x"8C660110",
x"C7E1021C",
x"8CC3FFEC",
x"C4600000",
x"44201801",
x"C7E10218",
x"C460FFFC",
x"44202001",
x"C7E10214",
x"C460FFF8",
x"44201001",
x"A1230002",
x"03E31820",
x"8C6703CC",
x"8CC5FFFC",
x"48BC006A",
x"C4E00000",
x"44030001",
x"C4E1FFFC",
x"44010002",
x"C7E502D8",
x"44052802",
x"44A43000",
x"E8D00003",
x"44C02806",
x"08001F8C",
x"44C02807",
x"8CC5FFF0",
x"C4A6FFFC",
x"E8A60003",
x"20030000",
x"08001FA0",
x"C7E502D4",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"08001F98",
x"44C02807",
x"C4A6FFF8",
x"E8A60003",
x"20030000",
x"08001FA0",
x"C8300003",
x"20030001",
x"08001FA0",
x"20030000",
x"48600047",
x"C4E0FFF8",
x"44040001",
x"C4E1FFF4",
x"44010002",
x"C7E502DC",
x"44052802",
x"44A33000",
x"E8D00003",
x"44C02806",
x"08001FAC",
x"44C02807",
x"C4A60000",
x"E8A60003",
x"20030000",
x"08001FBF",
x"C7E502D4",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"08001FB7",
x"44C02807",
x"C4A6FFF8",
x"E8A60003",
x"20030000",
x"08001FBF",
x"C8300003",
x"20030001",
x"08001FBF",
x"20030000",
x"48600025",
x"C4E0FFF0",
x"44020801",
x"C4E0FFEC",
x"44202802",
x"C7E102DC",
x"44A10802",
x"44231000",
x"E8500003",
x"44400806",
x"08001FCB",
x"44400807",
x"C4A20000",
x"E8220003",
x"20030000",
x"08001FDE",
x"C7E102D8",
x"44A10802",
x"44241000",
x"E8500003",
x"44400806",
x"08001FD6",
x"44400807",
x"C4A2FFFC",
x"E8220003",
x"20030000",
x"08001FDE",
x"C8100003",
x"20030001",
x"08001FDE",
x"20030000",
x"48600003",
x"20030000",
x"08001FE3",
x"E7E50208",
x"20030003",
x"08001FE6",
x"E7E00208",
x"20030002",
x"08001FE9",
x"E7E00208",
x"20030001",
x"0800203D",
x"20030002",
x"48A30010",
x"C4E00000",
x"E8100003",
x"20030000",
x"08001FFA",
x"C4E0FFFC",
x"44030802",
x"C4E0FFF8",
x"44040002",
x"44200800",
x"C4E0FFF4",
x"44020002",
x"44200000",
x"E7E00208",
x"20030001",
x"0800203D",
x"C4E00000",
x"C8100040",
x"C4E1FFFC",
x"44232802",
x"C4E1FFF8",
x"44240802",
x"44A12800",
x"C4E1FFF4",
x"44220802",
x"44A10800",
x"44633002",
x"8CC3FFF0",
x"C4650000",
x"44C53802",
x"44843002",
x"C465FFFC",
x"44C52802",
x"44E53800",
x"44423002",
x"C465FFF8",
x"44C52802",
x"44E53000",
x"8CC3FFF4",
x"48600003",
x"44C02806",
x"08002022",
x"44823802",
x"8CC3FFDC",
x"C4650000",
x"44E52802",
x"44C53000",
x"44432802",
x"C462FFFC",
x"44A21002",
x"44C23000",
x"44641802",
x"C462FFF8",
x"44622802",
x"44C52800",
x"20030003",
x"48A30003",
x"44B11001",
x"08002027",
x"44A01006",
x"44211802",
x"44020002",
x"44600001",
x"EA000003",
x"20030000",
x"0800203B",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"0800203A",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"0800203D",
x"20030000",
x"C7E00208",
x"48600003",
x"20030000",
x"08002047",
x"2003009C",
x"C4610000",
x"E8010003",
x"20030000",
x"08002047",
x"20030001",
x"4860000A",
x"A1230002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600003",
x"20030000",
x"E0000000",
x"21080001",
x"08001F6A",
x"20030098",
x"C4610000",
x"44010000",
x"C7E10134",
x"44201002",
x"C7E1021C",
x"44412800",
x"C7E10130",
x"44201002",
x"C7E10218",
x"44412000",
x"C7E1012C",
x"44200802",
x"C7E00214",
x"44201800",
x"8C850000",
x"AC240000",
x"48BD0003",
x"20030001",
x"080020DB",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08002075",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"0800208B",
x"E8500003",
x"44400006",
x"0800207E",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"0800208B",
x"E8300003",
x"44200006",
x"08002086",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"0800208B",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08002091",
x"20030000",
x"08002093",
x"8CC3FFE8",
x"080020D4",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080020A4",
x"20050001",
x"48650003",
x"20030001",
x"080020A8",
x"20030000",
x"080020D4",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"080020C6",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"080020CB",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080020D0",
x"20050001",
x"48650003",
x"20030001",
x"080020D4",
x"20030000",
x"48600006",
x"20050001",
x"40210008",
x"C0001E79",
x"20210008",
x"080020DB",
x"20030000",
x"48600004",
x"21080001",
x"8C240000",
x"08001F6A",
x"20030001",
x"E0000000",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600073",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600063",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600053",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600043",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600033",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600023",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600013",
x"216B0001",
x"A1630002",
x"4D432000",
x"489D0003",
x"20030000",
x"E0000000",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210004",
x"C0001F6A",
x"20210004",
x"48600003",
x"216B0001",
x"080020E1",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"20030001",
x"E0000000",
x"A1830002",
x"4DA35000",
x"8D440000",
x"489D0003",
x"20030000",
x"E0000000",
x"20030063",
x"AC2A0000",
x"48830003",
x"20030001",
x"080022AE",
x"A0830002",
x"03E31820",
x"8C650110",
x"C7E1021C",
x"8CA3FFEC",
x"C4600000",
x"44201801",
x"C7E10218",
x"C460FFFC",
x"44202001",
x"C7E10214",
x"C460FFF8",
x"44200801",
x"A0830002",
x"03E31820",
x"8C6603CC",
x"8CA4FFFC",
x"489C006A",
x"C4C00000",
x"44031001",
x"C4C0FFFC",
x"44403002",
x"C7E202D8",
x"44C21002",
x"44442800",
x"E8B00003",
x"44A01006",
x"0800218A",
x"44A01007",
x"8CA4FFF0",
x"C485FFFC",
x"E8450003",
x"20030000",
x"0800219E",
x"C7E202D4",
x"44C21002",
x"44412800",
x"E8B00003",
x"44A01006",
x"08002196",
x"44A01007",
x"C485FFF8",
x"E8450003",
x"20030000",
x"0800219E",
x"C8100003",
x"20030001",
x"0800219E",
x"20030000",
x"48600047",
x"C4C0FFF8",
x"44040001",
x"C4C6FFF4",
x"44062802",
x"C7E002DC",
x"44A00002",
x"44031000",
x"E8500003",
x"44400006",
x"080021AA",
x"44400007",
x"C4820000",
x"E8020003",
x"20030000",
x"080021BD",
x"C7E002D4",
x"44A00002",
x"44011000",
x"E8500003",
x"44400006",
x"080021B5",
x"44400007",
x"C482FFF8",
x"E8020003",
x"20030000",
x"080021BD",
x"C8D00003",
x"20030001",
x"080021BD",
x"20030000",
x"48600025",
x"C4C0FFF0",
x"44010001",
x"C4C5FFEC",
x"44051002",
x"C7E002DC",
x"44400002",
x"44030800",
x"E8300003",
x"44200006",
x"080021C9",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"080021DC",
x"C7E002D8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"080021D4",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"080021DC",
x"C8B00003",
x"20030001",
x"080021DC",
x"20030000",
x"48600003",
x"20030000",
x"080021E1",
x"E7E20208",
x"20030003",
x"080021E4",
x"E7E50208",
x"20030002",
x"080021E7",
x"E7E60208",
x"20030001",
x"0800223B",
x"20030002",
x"48830010",
x"C4C00000",
x"E8100003",
x"20030000",
x"080021F8",
x"C4C0FFFC",
x"44031002",
x"C4C0FFF8",
x"44040002",
x"44401000",
x"C4C0FFF4",
x"44010002",
x"44400000",
x"E7E00208",
x"20030001",
x"0800223B",
x"C4C00000",
x"C8100040",
x"C4C2FFFC",
x"44432802",
x"C4C2FFF8",
x"44441002",
x"44A22800",
x"C4C2FFF4",
x"44411002",
x"44A21000",
x"44633002",
x"8CA3FFF0",
x"C4650000",
x"44C53802",
x"44843002",
x"C465FFFC",
x"44C52802",
x"44E53800",
x"44213002",
x"C465FFF8",
x"44C52802",
x"44E53000",
x"8CA3FFF4",
x"48600003",
x"44C02806",
x"08002220",
x"44813802",
x"8CA3FFDC",
x"C4650000",
x"44E52802",
x"44C53000",
x"44232802",
x"C461FFFC",
x"44A10802",
x"44C13000",
x"44641802",
x"C461FFF8",
x"44612802",
x"44C52800",
x"20030003",
x"48830003",
x"44B10801",
x"08002225",
x"44A00806",
x"44421802",
x"44010002",
x"44600001",
x"EA000003",
x"20030000",
x"08002239",
x"8CA3FFE8",
x"48600007",
x"44000004",
x"44400801",
x"C4C0FFF0",
x"44200002",
x"E7E00208",
x"08002238",
x"44000004",
x"44400800",
x"C4C0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"0800223B",
x"20030000",
x"48600003",
x"20030000",
x"080022AE",
x"C7E10208",
x"20030094",
x"C4600000",
x"E8200003",
x"20030000",
x"080022AE",
x"8D44FFFC",
x"489D0003",
x"20030000",
x"080022AA",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860005A",
x"8D44FFF8",
x"489D0003",
x"20030000",
x"080022A8",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860004C",
x"8D44FFF4",
x"489D0003",
x"20030000",
x"080022A6",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860003E",
x"8D44FFF0",
x"489D0003",
x"20030000",
x"080022A4",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600030",
x"8D44FFEC",
x"489D0003",
x"20030000",
x"080022A2",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600022",
x"8D44FFE8",
x"489D0003",
x"20030000",
x"080022A0",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600014",
x"8D44FFE4",
x"489D0003",
x"20030000",
x"0800229E",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600006",
x"200B0008",
x"40210008",
x"C00020E1",
x"20210008",
x"0800229E",
x"20030001",
x"080022A0",
x"20030001",
x"080022A2",
x"20030001",
x"080022A4",
x"20030001",
x"080022A6",
x"20030001",
x"080022A8",
x"20030001",
x"080022AA",
x"20030001",
x"48600003",
x"20030000",
x"080022AE",
x"20030001",
x"48600003",
x"218C0001",
x"08002162",
x"8C2A0000",
x"8D44FFFC",
x"489D0003",
x"20030000",
x"08002318",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860005A",
x"8D44FFF8",
x"489D0003",
x"20030000",
x"08002316",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860004C",
x"8D44FFF4",
x"489D0003",
x"20030000",
x"08002314",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"4860003E",
x"8D44FFF0",
x"489D0003",
x"20030000",
x"08002312",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600030",
x"8D44FFEC",
x"489D0003",
x"20030000",
x"08002310",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600022",
x"8D44FFE8",
x"489D0003",
x"20030000",
x"0800230E",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600014",
x"8D44FFE4",
x"489D0003",
x"20030000",
x"0800230C",
x"A0830002",
x"03E31820",
x"8C640200",
x"20080000",
x"40210008",
x"C0001F6A",
x"20210008",
x"48600006",
x"200B0008",
x"40210008",
x"C00020E1",
x"20210008",
x"0800230C",
x"20030001",
x"0800230E",
x"20030001",
x"08002310",
x"20030001",
x"08002312",
x"20030001",
x"08002314",
x"20030001",
x"08002316",
x"20030001",
x"08002318",
x"20030001",
x"48600003",
x"218C0001",
x"08002162",
x"20030001",
x"E0000000",
x"A1630002",
x"4C835000",
x"495D0002",
x"E0000000",
x"A1430002",
x"03E31820",
x"8C670110",
x"C7E10270",
x"8CE3FFEC",
x"C4600000",
x"44203001",
x"C7E1026C",
x"C460FFFC",
x"44203801",
x"C7E10268",
x"C460FFF8",
x"44202801",
x"8CE3FFFC",
x"487C0087",
x"C5220000",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"08002338",
x"20060001",
x"C4A10000",
x"48660003",
x"44200007",
x"0800233D",
x"44200006",
x"44060001",
x"44021003",
x"C520FFFC",
x"44400002",
x"44070800",
x"E8300003",
x"44200006",
x"08002346",
x"44200007",
x"C4A1FFFC",
x"E8010003",
x"20080000",
x"08002357",
x"C520FFF8",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08002351",
x"44200007",
x"C4A1FFF8",
x"E8010003",
x"20080000",
x"08002357",
x"E7E20208",
x"20080001",
x"08002359",
x"20080000",
x"4900005B",
x"C522FFFC",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"08002362",
x"20060001",
x"C4A1FFFC",
x"48660003",
x"44200007",
x"08002367",
x"44200006",
x"44070001",
x"44021003",
x"C520FFF8",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08002370",
x"44200007",
x"C4A1FFF8",
x"E8010003",
x"20080000",
x"08002381",
x"C5200000",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"0800237B",
x"44200007",
x"C4A10000",
x"E8010003",
x"20080000",
x"08002381",
x"E7E20208",
x"20080001",
x"08002383",
x"20080000",
x"4900002F",
x"C522FFF8",
x"C8500027",
x"8CE5FFF0",
x"8CE3FFE8",
x"E8500003",
x"20060000",
x"0800238C",
x"20060001",
x"C4A1FFF8",
x"48660003",
x"44200007",
x"08002391",
x"44200006",
x"44050001",
x"44021003",
x"C5200000",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"0800239A",
x"44200007",
x"C4A10000",
x"E8010003",
x"20080000",
x"080023AB",
x"C520FFFC",
x"44400002",
x"44070800",
x"E8300003",
x"44200006",
x"080023A5",
x"44200007",
x"C4A1FFFC",
x"E8010003",
x"20080000",
x"080023AB",
x"E7E20208",
x"20080001",
x"080023AD",
x"20080000",
x"49000003",
x"20080000",
x"080023B1",
x"20080003",
x"080023B3",
x"20080002",
x"080023B5",
x"20080001",
x"08002440",
x"20080002",
x"4868001A",
x"8CE3FFF0",
x"C5200000",
x"C4640000",
x"44040802",
x"C520FFFC",
x"C463FFFC",
x"44030002",
x"44201000",
x"C520FFF8",
x"C461FFF8",
x"44010002",
x"44400000",
x"EA000003",
x"20080000",
x"080023D0",
x"44862002",
x"44671002",
x"44821000",
x"44250802",
x"44410800",
x"44200807",
x"44200003",
x"E7E00208",
x"20080001",
x"08002440",
x"C5210000",
x"C522FFFC",
x"C520FFF8",
x"44211802",
x"8CE5FFF0",
x"C4AA0000",
x"446A2002",
x"44421802",
x"C4ACFFFC",
x"446C1802",
x"44832000",
x"44001802",
x"C4ABFFF8",
x"446B1802",
x"44831800",
x"8CE6FFF4",
x"48C00003",
x"44604806",
x"080023F1",
x"44404002",
x"8CE5FFDC",
x"C4A40000",
x"45042002",
x"44644000",
x"44012002",
x"C4A3FFFC",
x"44831802",
x"45034000",
x"44222002",
x"C4A3FFF8",
x"44834802",
x"45094800",
x"C930004E",
x"44261802",
x"446A2002",
x"44471802",
x"446C1802",
x"44832000",
x"44051802",
x"446B1802",
x"44834000",
x"48C00003",
x"45001806",
x"08002411",
x"44072002",
x"44451802",
x"44832000",
x"8CE5FFDC",
x"C4A30000",
x"44832002",
x"44251802",
x"44060002",
x"44601800",
x"C4A0FFFC",
x"44600002",
x"44800000",
x"44271802",
x"44460802",
x"44611000",
x"C4A1FFF8",
x"44410802",
x"44010000",
x"44151802",
x"45031800",
x"44C60002",
x"440A0802",
x"44E70002",
x"440C0002",
x"44200800",
x"44A50002",
x"440B0002",
x"44200800",
x"48C00003",
x"44200006",
x"08002429",
x"44E51002",
x"8CE5FFDC",
x"C4A00000",
x"44400002",
x"44201000",
x"44A60802",
x"C4A0FFFC",
x"44200002",
x"44401000",
x"44C70802",
x"C4A0FFF8",
x"44200002",
x"44400000",
x"20050003",
x"48650003",
x"44110801",
x"0800242E",
x"44000806",
x"44631002",
x"45210002",
x"44400001",
x"EA000003",
x"20080000",
x"0800243E",
x"44000004",
x"8CE3FFE8",
x"48600003",
x"44000807",
x"0800243A",
x"44000806",
x"44230001",
x"44090003",
x"E7E00208",
x"20080001",
x"08002440",
x"20080000",
x"49000009",
x"A1430002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600002",
x"E0000000",
x"216B0001",
x"0800231D",
x"C7E00208",
x"AC240000",
x"EA000002",
x"080024E7",
x"C7E10210",
x"E8010002",
x"080024E7",
x"20030098",
x"C4610000",
x"44014800",
x"C5200000",
x"44090802",
x"C7E00270",
x"44202800",
x"C520FFFC",
x"44090802",
x"C7E0026C",
x"44202000",
x"C520FFF8",
x"44090802",
x"C7E00268",
x"44201800",
x"8C850000",
x"E4230004",
x"E4240008",
x"E425000C",
x"48BD0003",
x"20030001",
x"080024DC",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08002476",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"0800248C",
x"E8500003",
x"44400006",
x"0800247F",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"0800248C",
x"E8300003",
x"44200006",
x"08002487",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"0800248C",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"08002492",
x"20030000",
x"08002494",
x"8CC3FFE8",
x"080024D5",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080024A5",
x"20050001",
x"48650003",
x"20030001",
x"080024A9",
x"20030000",
x"080024D5",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"080024C7",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"080024CC",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"080024D1",
x"20050001",
x"48650003",
x"20030001",
x"080024D5",
x"20030000",
x"48600006",
x"20050001",
x"40210014",
x"C0001E79",
x"20210014",
x"080024DC",
x"20030000",
x"48600002",
x"080024E7",
x"E7E90210",
x"C425000C",
x"E7E5021C",
x"C4240008",
x"E7E40218",
x"C4230004",
x"E7E30214",
x"AFEA0220",
x"AFE8020C",
x"216B0001",
x"8C240000",
x"0800231D",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"AC290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"A1A30002",
x"4D831800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"21AD0001",
x"8C290000",
x"080024EA",
x"A1C30002",
x"4DE36000",
x"8D830000",
x"487D0002",
x"E0000000",
x"20040063",
x"AC290000",
x"48640053",
x"8D83FFFC",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF8",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF4",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF0",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFEC",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFE8",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFE4",
x"487D0002",
x"080025AD",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"200D0008",
x"8C290000",
x"40210008",
x"C00024EA",
x"20210008",
x"08002724",
x"A0630002",
x"03E31820",
x"8C660110",
x"C7E10270",
x"8CC3FFEC",
x"C4600000",
x"44202801",
x"C7E1026C",
x"C460FFFC",
x"44203001",
x"C7E10268",
x"C460FFF8",
x"44202001",
x"8CC4FFFC",
x"489C0087",
x"C5220000",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"080025C5",
x"20050001",
x"C4810000",
x"48650003",
x"44200007",
x"080025CA",
x"44200006",
x"44050001",
x"44021003",
x"C520FFFC",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"080025D3",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"080025E4",
x"C520FFF8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"080025DE",
x"44200007",
x"C481FFF8",
x"E8010003",
x"20030000",
x"080025E4",
x"E7E20208",
x"20030001",
x"080025E6",
x"20030000",
x"4860005B",
x"C522FFFC",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"080025EF",
x"20050001",
x"C481FFFC",
x"48650003",
x"44200007",
x"080025F4",
x"44200006",
x"44060001",
x"44021003",
x"C520FFF8",
x"44400002",
x"44040800",
x"E8300003",
x"44200006",
x"080025FD",
x"44200007",
x"C481FFF8",
x"E8010003",
x"20030000",
x"0800260E",
x"C5200000",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08002608",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"0800260E",
x"E7E20208",
x"20030001",
x"08002610",
x"20030000",
x"4860002F",
x"C522FFF8",
x"C8500027",
x"8CC4FFF0",
x"8CC3FFE8",
x"E8500003",
x"20050000",
x"08002619",
x"20050001",
x"C481FFF8",
x"48650003",
x"44200007",
x"0800261E",
x"44200006",
x"44040001",
x"44021003",
x"C5200000",
x"44400002",
x"44050800",
x"E8300003",
x"44200006",
x"08002627",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"08002638",
x"C520FFFC",
x"44400002",
x"44060800",
x"E8300003",
x"44200006",
x"08002632",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"08002638",
x"E7E20208",
x"20030001",
x"0800263A",
x"20030000",
x"48600003",
x"20030000",
x"0800263E",
x"20030003",
x"08002640",
x"20030002",
x"08002642",
x"20030001",
x"080026CD",
x"20030002",
x"4883001A",
x"8CC3FFF0",
x"C5200000",
x"C4670000",
x"44070802",
x"C520FFFC",
x"C463FFFC",
x"44030002",
x"44201000",
x"C520FFF8",
x"C461FFF8",
x"44010002",
x"44400000",
x"EA000003",
x"20030000",
x"0800265D",
x"44E52802",
x"44661002",
x"44A21000",
x"44240802",
x"44410800",
x"44200807",
x"44200003",
x"E7E00208",
x"20030001",
x"080026CD",
x"C5210000",
x"C522FFFC",
x"C520FFF8",
x"44211802",
x"8CC3FFF0",
x"C4690000",
x"44693802",
x"44421802",
x"C46BFFFC",
x"446B1802",
x"44E33800",
x"44001802",
x"C46AFFF8",
x"446A1802",
x"44E31800",
x"8CC5FFF4",
x"48A00003",
x"44604006",
x"0800267E",
x"44404002",
x"8CC3FFDC",
x"C4670000",
x"45073802",
x"44674000",
x"44013802",
x"C463FFFC",
x"44E31802",
x"45036000",
x"44223802",
x"C463FFF8",
x"44E34002",
x"45884000",
x"C910004E",
x"44251802",
x"44693802",
x"44461802",
x"446B1802",
x"44E33800",
x"44041802",
x"446A1802",
x"44E33800",
x"48A00003",
x"44E01806",
x"0800269E",
x"44066002",
x"44441802",
x"45836000",
x"8CC3FFDC",
x"C4630000",
x"45831802",
x"44246002",
x"44050002",
x"45806000",
x"C460FFFC",
x"45800002",
x"44600000",
x"44261802",
x"44450802",
x"44611000",
x"C461FFF8",
x"44410802",
x"44010000",
x"44151802",
x"44E31800",
x"44A50002",
x"44090802",
x"44C60002",
x"440B0002",
x"44200800",
x"44840002",
x"440A0002",
x"44200800",
x"48A00003",
x"44200006",
x"080026B6",
x"44C41002",
x"8CC3FFDC",
x"C4600000",
x"44400002",
x"44201000",
x"44850802",
x"C460FFFC",
x"44200002",
x"44401000",
x"44A60802",
x"C460FFF8",
x"44200002",
x"44400000",
x"20030003",
x"48830003",
x"44110801",
x"080026BB",
x"44000806",
x"44631002",
x"45010002",
x"44400001",
x"EA000003",
x"20030000",
x"080026CB",
x"44000004",
x"8CC3FFE8",
x"48600003",
x"44000807",
x"080026C7",
x"44000806",
x"44230001",
x"44080003",
x"E7E00208",
x"20030001",
x"080026CD",
x"20030000",
x"48600002",
x"08002724",
x"C7E00208",
x"C7E10210",
x"E8010002",
x"08002724",
x"8D83FFFC",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF8",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF4",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFF0",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFEC",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFE8",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"8D83FFE4",
x"487D0002",
x"08002724",
x"A0630002",
x"03E31820",
x"8C640200",
x"200B0000",
x"8C290000",
x"40210008",
x"C000231D",
x"20210008",
x"200D0008",
x"8C290000",
x"40210008",
x"C00024EA",
x"20210008",
x"21CE0001",
x"8C290000",
x"08002554",
x"A1430002",
x"4C834800",
x"493D0002",
x"E0000000",
x"A1230002",
x"03E31820",
x"8C660110",
x"8CC5FFD8",
x"C4A30000",
x"C4A4FFFC",
x"C4A2FFF8",
x"A1230002",
x"4D633800",
x"8CC3FFFC",
x"487C006A",
x"C4E00000",
x"44030001",
x"C4E1FFFC",
x"44010002",
x"C585FFFC",
x"44052802",
x"44A43000",
x"E8D00003",
x"44C02806",
x"08002741",
x"44C02807",
x"8CC3FFF0",
x"C466FFFC",
x"E8A60003",
x"20080000",
x"08002755",
x"C585FFF8",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"0800274D",
x"44C02807",
x"C466FFF8",
x"E8A60003",
x"20080000",
x"08002755",
x"C8300003",
x"20080001",
x"08002755",
x"20080000",
x"49000047",
x"C4E0FFF8",
x"44040001",
x"C4E1FFF4",
x"44010002",
x"C5850000",
x"44052802",
x"44A33000",
x"E8D00003",
x"44C02806",
x"08002761",
x"44C02807",
x"C4660000",
x"E8A60003",
x"20080000",
x"08002774",
x"C585FFF8",
x"44052802",
x"44A23000",
x"E8D00003",
x"44C02806",
x"0800276C",
x"44C02807",
x"C466FFF8",
x"E8A60003",
x"20080000",
x"08002774",
x"C8300003",
x"20080001",
x"08002774",
x"20080000",
x"49000025",
x"C4E0FFF0",
x"44020801",
x"C4E0FFEC",
x"44202802",
x"C5810000",
x"44A10802",
x"44231000",
x"E8500003",
x"44400806",
x"08002780",
x"44400807",
x"C4620000",
x"E8220003",
x"20080000",
x"08002793",
x"C581FFFC",
x"44A10802",
x"44241000",
x"E8500003",
x"44400806",
x"0800278B",
x"44400807",
x"C462FFFC",
x"E8220003",
x"20080000",
x"08002793",
x"C8100003",
x"20080001",
x"08002793",
x"20080000",
x"49000003",
x"20080000",
x"08002798",
x"E7E50208",
x"20080003",
x"0800279B",
x"E7E00208",
x"20080002",
x"0800279E",
x"E7E00208",
x"20080001",
x"080027CB",
x"20080002",
x"4868000A",
x"C4E10000",
x"E8300003",
x"20080000",
x"080027A9",
x"C4A0FFF4",
x"44200002",
x"E7E00208",
x"20080001",
x"080027CB",
x"C4E50000",
x"C8B0001F",
x"C4E0FFFC",
x"44030802",
x"C4E0FFF8",
x"44040002",
x"44200800",
x"C4E0FFF4",
x"44020002",
x"44200800",
x"C4A0FFF4",
x"44211002",
x"44A00002",
x"44400001",
x"EA000003",
x"20080000",
x"080027C9",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"080027C8",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20080001",
x"080027CB",
x"20080000",
x"49000009",
x"A1230002",
x"03E31820",
x"8C630110",
x"8C63FFE8",
x"48600002",
x"E0000000",
x"214A0001",
x"08002727",
x"C7E00208",
x"AC240000",
x"EA000002",
x"08002872",
x"C7E10210",
x"E8010002",
x"08002872",
x"20030098",
x"C4610000",
x"44014800",
x"C5800000",
x"44090802",
x"C7E0027C",
x"44202800",
x"C580FFFC",
x"44090802",
x"C7E00278",
x"44202000",
x"C580FFF8",
x"44090802",
x"C7E00274",
x"44201800",
x"8C850000",
x"E4230004",
x"E4240008",
x"E425000C",
x"48BD0003",
x"20030001",
x"08002867",
x"A0A30002",
x"03E31820",
x"8C660110",
x"8CC3FFEC",
x"C4600000",
x"44A00001",
x"C461FFFC",
x"44811001",
x"C461FFF8",
x"44610801",
x"8CC5FFFC",
x"48BC0024",
x"E8100003",
x"44003006",
x"08002801",
x"44003007",
x"8CC3FFF0",
x"C4600000",
x"E8C00003",
x"20050000",
x"08002817",
x"E8500003",
x"44400006",
x"0800280A",
x"44400007",
x"C462FFFC",
x"E8020003",
x"20050000",
x"08002817",
x"E8300003",
x"44200006",
x"08002812",
x"44200007",
x"C461FFF8",
x"E8010003",
x"20050000",
x"08002817",
x"20050001",
x"48A00007",
x"8CC3FFE8",
x"48600003",
x"20030001",
x"0800281D",
x"20030000",
x"0800281F",
x"8CC3FFE8",
x"08002860",
x"20030002",
x"48A30014",
x"8CC3FFF0",
x"C4660000",
x"44C03002",
x"C460FFFC",
x"44020002",
x"44C01000",
x"C460FFF8",
x"44010002",
x"44400000",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"08002830",
x"20050001",
x"48650003",
x"20030001",
x"08002834",
x"20030000",
x"08002860",
x"44003802",
x"8CC3FFF0",
x"C4660000",
x"44E64002",
x"44423802",
x"C466FFFC",
x"44E63002",
x"45064000",
x"44213802",
x"C466FFF8",
x"44E63002",
x"45063800",
x"8CC3FFF4",
x"48600003",
x"44E03006",
x"08002852",
x"44414002",
x"8CC3FFDC",
x"C4660000",
x"45063002",
x"44E63800",
x"44203002",
x"C461FFFC",
x"44C10802",
x"44E13800",
x"44020802",
x"C460FFF8",
x"44203002",
x"44E63000",
x"20030003",
x"48A30003",
x"44D10001",
x"08002857",
x"44C00006",
x"8CC3FFE8",
x"E8100003",
x"20050000",
x"0800285C",
x"20050001",
x"48650003",
x"20030001",
x"08002860",
x"20030000",
x"48600006",
x"20050001",
x"40210014",
x"C0001E79",
x"20210014",
x"08002867",
x"20030000",
x"48600002",
x"08002872",
x"E7E90210",
x"C425000C",
x"E7E5021C",
x"C4240008",
x"E7E40218",
x"C4230004",
x"E7E30214",
x"AFE90220",
x"AFE8020C",
x"214A0001",
x"8C240000",
x"08002727",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"A2030002",
x"4DE31800",
x"487D0002",
x"E0000000",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"21AB0000",
x"21CC0000",
x"40210004",
x"C0002727",
x"20210004",
x"22100001",
x"08002875",
x"A2630002",
x"4E837800",
x"8DE30000",
x"487D0002",
x"E0000000",
x"20040063",
x"4864005A",
x"8DE3FFFC",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF8",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF4",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF0",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFEC",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFE8",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFE4",
x"487D0002",
x"08002945",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20100008",
x"222D0000",
x"224E0000",
x"C0002875",
x"20210004",
x"08002A44",
x"A0640002",
x"03E42020",
x"8C860110",
x"8CC5FFD8",
x"C4A20000",
x"C4A3FFFC",
x"C4A1FFF8",
x"A0630002",
x"4E233800",
x"8CC4FFFC",
x"489C006A",
x"C4E00000",
x"44022001",
x"C4E0FFFC",
x"44803002",
x"C644FFFC",
x"44C42002",
x"44832800",
x"E8B00003",
x"44A02006",
x"0800295C",
x"44A02007",
x"8CC4FFF0",
x"C485FFFC",
x"E8850003",
x"20030000",
x"08002970",
x"C644FFF8",
x"44C42002",
x"44812800",
x"E8B00003",
x"44A02006",
x"08002968",
x"44A02007",
x"C485FFF8",
x"E8850003",
x"20030000",
x"08002970",
x"C8100003",
x"20030001",
x"08002970",
x"20030000",
x"48600047",
x"C4E0FFF8",
x"44030001",
x"C4E6FFF4",
x"44062802",
x"C6400000",
x"44A00002",
x"44022000",
x"E8900003",
x"44800006",
x"0800297C",
x"44800007",
x"C4840000",
x"E8040003",
x"20030000",
x"0800298F",
x"C640FFF8",
x"44A00002",
x"44012000",
x"E8900003",
x"44800006",
x"08002987",
x"44800007",
x"C484FFF8",
x"E8040003",
x"20030000",
x"0800298F",
x"C8D00003",
x"20030001",
x"0800298F",
x"20030000",
x"48600025",
x"C4E0FFF0",
x"44010001",
x"C4E5FFEC",
x"44052002",
x"C6400000",
x"44800002",
x"44020800",
x"E8300003",
x"44200006",
x"0800299B",
x"44200007",
x"C4810000",
x"E8010003",
x"20030000",
x"080029AE",
x"C640FFFC",
x"44800002",
x"44030800",
x"E8300003",
x"44200006",
x"080029A6",
x"44200007",
x"C481FFFC",
x"E8010003",
x"20030000",
x"080029AE",
x"C8B00003",
x"20030001",
x"080029AE",
x"20030000",
x"48600003",
x"20030000",
x"080029B3",
x"E7E40208",
x"20030003",
x"080029B6",
x"E7E50208",
x"20030002",
x"080029B9",
x"E7E60208",
x"20030001",
x"080029E6",
x"20030002",
x"4883000A",
x"C4E10000",
x"E8300003",
x"20030000",
x"080029C4",
x"C4A0FFF4",
x"44200002",
x"E7E00208",
x"20030001",
x"080029E6",
x"C4E40000",
x"C890001F",
x"C4E0FFFC",
x"44021002",
x"C4E0FFF8",
x"44030002",
x"44401000",
x"C4E0FFF4",
x"44010002",
x"44400800",
x"C4A0FFF4",
x"44211002",
x"44800002",
x"44400001",
x"EA000003",
x"20030000",
x"080029E4",
x"8CC3FFE8",
x"48600007",
x"44000004",
x"44200801",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"080029E3",
x"44000004",
x"44200800",
x"C4E0FFF0",
x"44200002",
x"E7E00208",
x"20030001",
x"080029E6",
x"20030000",
x"48600002",
x"08002A44",
x"C7E00208",
x"C7E10210",
x"E8010002",
x"08002A44",
x"8DE3FFFC",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF8",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF4",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFF0",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFEC",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFE8",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20210004",
x"8DE3FFE4",
x"487D0002",
x"08002A44",
x"A0630002",
x"03E31820",
x"8C640200",
x"200A0000",
x"222B0000",
x"224C0000",
x"40210004",
x"C0002727",
x"20100008",
x"222D0000",
x"224E0000",
x"C0002875",
x"20210004",
x"22730001",
x"080028E6",
x"6AA00064",
x"A2A30002",
x"03E31820",
x"8C7706B4",
x"8EF8FFFC",
x"200300D4",
x"C4600000",
x"E7E00210",
x"20130000",
x"8FF40204",
x"8F11FFFC",
x"8F120000",
x"40210004",
x"C00028E6",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"08002A61",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"08002A61",
x"20030001",
x"48600002",
x"08002AA8",
x"8FE30220",
x"A0640002",
x"8FE3020C",
x"00831820",
x"8EE40000",
x"48640040",
x"200C0000",
x"8FED0204",
x"40210004",
x"C0002162",
x"20210004",
x"48600039",
x"8F030000",
x"C7E0022C",
x"C4620000",
x"44020802",
x"C7E00228",
x"C464FFFC",
x"44040002",
x"44200800",
x"C7E00224",
x"C463FFF8",
x"44030002",
x"44200800",
x"C6E0FFF8",
x"440B2802",
x"44A10802",
x"C6C50000",
x"44A22802",
x"C6C2FFFC",
x"44441002",
x"44A22000",
x"C6C2FFF8",
x"44431002",
x"44821000",
x"44020002",
x"EA010002",
x"08002A98",
x"C7E30250",
x"C7E20238",
x"44221002",
x"44621000",
x"E7E20250",
x"C7E3024C",
x"C7E20234",
x"44221002",
x"44621000",
x"E7E2024C",
x"C7E30248",
x"C7E20230",
x"44220802",
x"44610800",
x"E7E10248",
x"EA000002",
x"08002AA6",
x"44000002",
x"44000002",
x"440A0002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"08002AA7",
x"08002AA8",
x"42B50001",
x"08002A46",
x"E0000000",
x"20030004",
x"68790415",
x"200300D4",
x"C4600000",
x"E7E00210",
x"200E0000",
x"8FEF0204",
x"22C90000",
x"40210004",
x"C0002554",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"08002AC2",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"08002AC2",
x"20030001",
x"48600023",
x"2004FFFF",
x"A3230002",
x"6E632000",
x"4B200002",
x"E0000000",
x"C6C10000",
x"C7E00134",
x"44201002",
x"C6C1FFFC",
x"C7E00130",
x"44200002",
x"44401000",
x"C6C1FFF8",
x"C7E0012C",
x"44200002",
x"44400000",
x"44000007",
x"EA000002",
x"E0000000",
x"44000802",
x"44200002",
x"440D0802",
x"C7E00138",
x"44200002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"E0000000",
x"8FE70220",
x"A0E30002",
x"03E31820",
x"8C630110",
x"8C7EFFF8",
x"8C7AFFE4",
x"C7400000",
x"440D5802",
x"8C64FFFC",
x"489C0016",
x"8FE4020C",
x"E7F0022C",
x"E7F00228",
x"E7F00224",
x"40850001",
x"A0A40002",
x"02C40831",
x"C8300008",
x"EA010004",
x"200400A0",
x"C4800000",
x"08002AFD",
x"200400C8",
x"C4800000",
x"08002AFF",
x"46000006",
x"44000007",
x"A0A40002",
x"03E42020",
x"E480022C",
x"08002B5B",
x"20050002",
x"4885000C",
x"8C64FFF0",
x"C4800000",
x"44000007",
x"E7E0022C",
x"C480FFFC",
x"44000007",
x"E7E00228",
x"C480FFF8",
x"44000007",
x"E7E00224",
x"08002B5B",
x"C7E1021C",
x"8C64FFEC",
x"C4800000",
x"44202001",
x"C7E10218",
x"C480FFFC",
x"44201801",
x"C7E10214",
x"C480FFF8",
x"44200001",
x"8C64FFF0",
x"C4810000",
x"44810802",
x"C482FFFC",
x"44622802",
x"C482FFF8",
x"44023802",
x"8C64FFF4",
x"48800005",
x"E7E1022C",
x"E7E50228",
x"E7E70224",
x"08002B41",
x"8C64FFDC",
x"C482FFF8",
x"44623002",
x"C482FFFC",
x"44021002",
x"44C21000",
x"44551002",
x"44220800",
x"E7E1022C",
x"C481FFF8",
x"44811002",
x"C4810000",
x"44010002",
x"44400000",
x"44150002",
x"44A00000",
x"E7E00228",
x"C480FFFC",
x"44800802",
x"C4800000",
x"44600002",
x"44200000",
x"44150002",
x"44E00000",
x"E7E00224",
x"8C64FFE8",
x"C7E2022C",
x"44420802",
x"C7E00228",
x"44000002",
x"44200800",
x"C7E00224",
x"44000002",
x"44200000",
x"44000804",
x"C8300006",
x"48800003",
x"46210003",
x"08002B50",
x"46810003",
x"08002B53",
x"200400C8",
x"C4800000",
x"44400802",
x"E7E1022C",
x"C7E10228",
x"44200802",
x"E7E10228",
x"C7E10224",
x"44200002",
x"E7E00224",
x"C7E0021C",
x"E7E00270",
x"C7E00218",
x"E7E0026C",
x"C7E00214",
x"E7E00268",
x"8C640000",
x"8C65FFE0",
x"C4A00000",
x"E7E00238",
x"C4A0FFFC",
x"E7E00234",
x"C4A0FFF8",
x"E7E00230",
x"489C0028",
x"C7E1021C",
x"8C65FFEC",
x"C4A00000",
x"44202801",
x"2003002C",
x"C4690000",
x"44A90002",
x"40210004",
x"C0000051",
x"20030028",
x"C4660000",
x"44060002",
x"44A04001",
x"20030034",
x"C4650000",
x"C7E10214",
x"C4A0FFF8",
x"44203801",
x"44E90002",
x"C0000051",
x"20210004",
x"44060002",
x"44E00801",
x"E9050008",
x"E8250004",
x"200300D8",
x"C4600000",
x"08002B88",
x"200300DC",
x"C4600000",
x"08002B8F",
x"E8250004",
x"200300DC",
x"C4600000",
x"08002B8F",
x"200300D8",
x"C4600000",
x"E7E00234",
x"08002DAB",
x"20050002",
x"48850082",
x"C7E10218",
x"20030030",
x"C4600000",
x"44201002",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"08002B9F",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08002BC5",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002BB6",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002BB1",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BB6",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BC5",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002BC0",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BC5",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BE8",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002BD9",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002BD4",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BD9",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BE8",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002BE3",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002BE8",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8600006",
x"EA020003",
x"20030000",
x"08002BED",
x"20030001",
x"08002BF2",
x"EA020003",
x"20030001",
x"08002BF2",
x"20030000",
x"E8600003",
x"44000806",
x"08002BF6",
x"47A00801",
x"EAC10003",
x"44200006",
x"08002BFA",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"08002C0D",
x"44000806",
x"44210002",
x"47600802",
x"E7E10238",
x"46200001",
x"47600002",
x"E7E00234",
x"08002DAB",
x"20050003",
x"48850095",
x"C7E1021C",
x"8C63FFEC",
x"C4600000",
x"44200001",
x"C7E20214",
x"C461FFF8",
x"44410801",
x"44000002",
x"44210802",
x"44010000",
x"44000004",
x"20030034",
x"C4610000",
x"44010003",
x"E4200000",
x"40210008",
x"C0000051",
x"20210008",
x"44000806",
x"C4200000",
x"44010001",
x"441E0002",
x"46C01001",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"08002C35",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08002C5B",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002C4C",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002C47",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C4C",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C5B",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002C56",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C5B",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C7E",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002C6F",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002C6A",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C6F",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C7E",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002C79",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08002C7E",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8600006",
x"EA020003",
x"20030000",
x"08002C83",
x"20030001",
x"08002C88",
x"EA020003",
x"20030001",
x"08002C88",
x"20030000",
x"E8600003",
x"44000806",
x"08002C8C",
x"47A00801",
x"EAC10003",
x"44200006",
x"08002C90",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"08002CA3",
x"44000806",
x"44210002",
x"441B0802",
x"E7E10234",
x"46200001",
x"441B0002",
x"E7E00230",
x"08002DAB",
x"20050004",
x"48850100",
x"C7E1021C",
x"8C66FFEC",
x"C4C00000",
x"44200801",
x"8C65FFF0",
x"C4A00000",
x"44000004",
x"44200802",
x"C7E20214",
x"C4C0FFF8",
x"44401001",
x"C4A0FFF8",
x"44000004",
x"44401002",
x"44211802",
x"44420002",
x"44602800",
x"E8300003",
x"44200006",
x"08002CC1",
x"44200007",
x"2003008C",
x"C4660000",
x"E806005D",
x"44410803",
x"E8300003",
x"44200006",
x"08002CC9",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"08002CCE",
x"2003FFFF",
x"08002CD0",
x"20030001",
x"48600003",
x"44001806",
x"08002CD4",
x"46201803",
x"44630002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44202002",
x"20040078",
x"C4810000",
x"44220800",
x"44811003",
x"20040074",
x"C4810000",
x"44202002",
x"20040070",
x"C4810000",
x"44220800",
x"44811003",
x"2004006C",
x"C4810000",
x"44202002",
x"20040068",
x"C4810000",
x"44220800",
x"44811003",
x"20040064",
x"C4810000",
x"44202002",
x"47820800",
x"44811003",
x"20040060",
x"C4810000",
x"44202002",
x"2004005C",
x"C4810000",
x"44220800",
x"44811003",
x"20040058",
x"C4810000",
x"44202002",
x"20040054",
x"C4810000",
x"44220800",
x"44811003",
x"20040050",
x"C4810000",
x"44202002",
x"47220800",
x"44810803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44202002",
x"47020800",
x"44810803",
x"46E10800",
x"44010003",
x"46200000",
x"44600803",
x"68030006",
x"68600003",
x"44200006",
x"08002D19",
x"47E10001",
x"08002D1B",
x"46C10001",
x"20030044",
x"C4610000",
x"44010002",
x"441E0003",
x"08002D22",
x"20030088",
x"C4600000",
x"E4200004",
x"4021000C",
x"C0000051",
x"2021000C",
x"44000806",
x"C4200004",
x"44013801",
x"C7E10218",
x"C4C0FFFC",
x"44200801",
x"C4A0FFFC",
x"44000004",
x"44200802",
x"E8B00003",
x"44A00006",
x"08002D33",
x"44A00007",
x"E806005D",
x"44250803",
x"E8300003",
x"44200006",
x"08002D39",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"08002D3E",
x"2003FFFF",
x"08002D40",
x"20030001",
x"48600003",
x"44002006",
x"08002D44",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44610803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800003",
x"68030006",
x"68600003",
x"44000806",
x"08002D89",
x"47E00801",
x"08002D8B",
x"46C00801",
x"20030044",
x"C4600000",
x"44200002",
x"441E0003",
x"08002D92",
x"20030088",
x"C4600000",
x"E4200008",
x"40210010",
x"C0000051",
x"20210010",
x"44000806",
x"C4200008",
x"44010001",
x"2003003C",
x"C4620000",
x"46A70801",
x"44210802",
x"44410801",
x"46A00001",
x"44000002",
x"44200801",
x"E8300003",
x"44200006",
x"08002DA5",
x"46000006",
x"47600802",
x"20030038",
x"C4600000",
x"44200003",
x"E7E00230",
x"08002DAB",
x"A0E40002",
x"8FE3020C",
x"00832020",
x"A3230002",
x"6E632000",
x"A3230002",
x"4E831800",
x"C7E0021C",
x"E4600000",
x"C7E00218",
x"E460FFFC",
x"C7E00214",
x"E460FFF8",
x"C7400000",
x"E8150023",
x"20040001",
x"A3230002",
x"6E432000",
x"A3230002",
x"4E231800",
x"C7E00238",
x"E4600000",
x"C7E00234",
x"E460FFFC",
x"C7E00230",
x"E460FFF8",
x"A3230002",
x"4E232000",
x"20030024",
x"C4600000",
x"440B0002",
x"C4810000",
x"44200802",
x"E4810000",
x"C481FFFC",
x"44200802",
x"E481FFFC",
x"C481FFF8",
x"44200002",
x"E480FFF8",
x"A3230002",
x"4E031800",
x"C7E0022C",
x"E4600000",
x"C7E00228",
x"E460FFFC",
x"C7E00224",
x"E460FFF8",
x"08002DDF",
x"20040000",
x"A3230002",
x"6E432000",
x"20030020",
x"C4630000",
x"C6C10000",
x"C7E0022C",
x"44202802",
x"C6C4FFFC",
x"C7E20228",
x"44821002",
x"44A22800",
x"C6C4FFF8",
x"C7E20224",
x"44821002",
x"44A21000",
x"44621002",
x"44400002",
x"44200000",
x"E6C00000",
x"C6C1FFFC",
x"C7E00228",
x"44400002",
x"44200000",
x"E6C0FFFC",
x"C6C1FFF8",
x"C7E00224",
x"44400002",
x"44200000",
x"E6C0FFF8",
x"C740FFFC",
x"45A05002",
x"200C0000",
x"8FED0204",
x"40210010",
x"C0002162",
x"20210010",
x"48600037",
x"C7E1022C",
x"C7E00134",
x"44201002",
x"C7E10228",
x"C7E30130",
x"44230802",
x"44412000",
x"C7E10224",
x"C7E2012C",
x"44220802",
x"44810800",
x"44200807",
x"442B0802",
x"C6C40000",
x"44802002",
x"C6C0FFFC",
x"44030002",
x"44801800",
x"C6C0FFF8",
x"44020002",
x"44600000",
x"44000007",
x"EA010002",
x"08002E29",
x"C7E30250",
x"C7E20238",
x"44221002",
x"44621000",
x"E7E20250",
x"C7E3024C",
x"C7E20234",
x"44221002",
x"44621000",
x"E7E2024C",
x"C7E30248",
x"C7E20230",
x"44220802",
x"44610800",
x"E7E10248",
x"EA000002",
x"08002E37",
x"44000002",
x"44000002",
x"440A0002",
x"C7E10250",
x"44200800",
x"E7E10250",
x"C7E1024C",
x"44200800",
x"E7E1024C",
x"C7E10248",
x"44200000",
x"E7E00248",
x"08002E38",
x"C7E0021C",
x"E7E0027C",
x"C7E00218",
x"E7E00278",
x"C7E00214",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7E1021C",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C7E10218",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C7E10214",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08002E8C",
x"20050002",
x"68A60002",
x"08002E8C",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"08002E86",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08002E8B",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"43E3021C",
x"40210010",
x"C0001DDC",
x"20210010",
x"08002E92",
x"8FE306B8",
x"40630001",
x"AC36000C",
x"AC300010",
x"AC350014",
x"AC370018",
x"AC31001C",
x"AC320020",
x"AC330024",
x"AC340028",
x"AC38002C",
x"AC330030",
x"20750000",
x"40210038",
x"C0002A46",
x"20210038",
x"200300A4",
x"C4600000",
x"E80D0002",
x"E0000000",
x"20030004",
x"6B230002",
x"08002EAE",
x"23230001",
x"2004FFFF",
x"A0630002",
x"8C330030",
x"6E632000",
x"20030002",
x"4BC30011",
x"C7400000",
x"46200001",
x"45A06802",
x"23390001",
x"C7E00210",
x"45C07000",
x"8C38002C",
x"8C340028",
x"8C330024",
x"8C320020",
x"8C31001C",
x"8C370018",
x"8C350014",
x"8C300010",
x"8C36000C",
x"08002AAB",
x"E0000000",
x"E0000000",
x"200400D4",
x"C4800000",
x"E7E00210",
x"20130000",
x"8FF40204",
x"20710000",
x"22B20000",
x"40210004",
x"C00028E6",
x"20210004",
x"C7E00210",
x"20030094",
x"C4610000",
x"E8200003",
x"20030000",
x"08002ED8",
x"20030090",
x"C4610000",
x"E8010003",
x"20030000",
x"08002ED8",
x"20030001",
x"48600002",
x"E0000000",
x"8FE30220",
x"A0630002",
x"03E31820",
x"8C6E0110",
x"8DC3FFFC",
x"487C0016",
x"8FE3020C",
x"E7F0022C",
x"E7F00228",
x"E7F00224",
x"40640001",
x"A0830002",
x"02A30831",
x"C8300008",
x"EA010004",
x"200300A0",
x"C4600000",
x"08002EEE",
x"200300C8",
x"C4600000",
x"08002EF0",
x"46000006",
x"44000007",
x"A0830002",
x"03E31820",
x"E460022C",
x"08002F4C",
x"20040002",
x"4864000C",
x"8DC3FFF0",
x"C4600000",
x"44000007",
x"E7E0022C",
x"C460FFFC",
x"44000007",
x"E7E00228",
x"C460FFF8",
x"44000007",
x"E7E00224",
x"08002F4C",
x"C7E1021C",
x"8DC3FFEC",
x"C4600000",
x"44202001",
x"C7E10218",
x"C460FFFC",
x"44201801",
x"C7E10214",
x"C460FFF8",
x"44200001",
x"8DC3FFF0",
x"C4610000",
x"44811002",
x"C461FFFC",
x"44613002",
x"C461FFF8",
x"44013802",
x"8DC3FFF4",
x"48600005",
x"E7E2022C",
x"E7E60228",
x"E7E70224",
x"08002F32",
x"8DC3FFDC",
x"C461FFF8",
x"44612802",
x"C461FFFC",
x"44010802",
x"44A10800",
x"44350802",
x"44410800",
x"E7E1022C",
x"C461FFF8",
x"44811002",
x"C4610000",
x"44010002",
x"44400000",
x"44150002",
x"44C00000",
x"E7E00228",
x"C460FFFC",
x"44800802",
x"C4600000",
x"44600002",
x"44200000",
x"44150002",
x"44E00000",
x"E7E00224",
x"8DC3FFE8",
x"C7E2022C",
x"44420802",
x"C7E00228",
x"44000002",
x"44200800",
x"C7E00224",
x"44000002",
x"44200000",
x"44000804",
x"C8300006",
x"48600003",
x"46210003",
x"08002F41",
x"46810003",
x"08002F44",
x"200300C8",
x"C4600000",
x"44400802",
x"E7E1022C",
x"C7E10228",
x"44200802",
x"E7E10228",
x"C7E10224",
x"44200002",
x"E7E00224",
x"8DC30000",
x"8DC4FFE0",
x"C4800000",
x"E7E00238",
x"C480FFFC",
x"E7E00234",
x"C480FFF8",
x"E7E00230",
x"487C0028",
x"C7E1021C",
x"8DC5FFEC",
x"C4A00000",
x"44202801",
x"2003002C",
x"C4690000",
x"44A90002",
x"40210004",
x"C0000051",
x"20030028",
x"C4680000",
x"44080002",
x"44A03801",
x"20030034",
x"C4660000",
x"C7E10214",
x"C4A0FFF8",
x"44202801",
x"44A90002",
x"C0000051",
x"20210004",
x"44080002",
x"44A00801",
x"E8E60008",
x"E8260004",
x"200300D8",
x"C4600000",
x"08002F73",
x"200300DC",
x"C4600000",
x"08002F7A",
x"E8260004",
x"200300DC",
x"C4600000",
x"08002F7A",
x"200300D8",
x"C4600000",
x"E7E00234",
x"08003196",
x"20040002",
x"48640082",
x"C7E10218",
x"20030030",
x"C4600000",
x"44201002",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"08002F8A",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08002FB0",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002FA1",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002F9C",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FA1",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FB0",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002FAB",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FB0",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FD3",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"08002FC4",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002FBF",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FC4",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FD3",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08002FCE",
x"443D0800",
x"40210004",
x"C0000DE4",
x"20210004",
x"08002FD3",
x"443D0801",
x"40210004",
x"C0000DE4",
x"20210004",
x"E8600006",
x"EA020003",
x"20030000",
x"08002FD8",
x"20030001",
x"08002FDD",
x"EA020003",
x"20030001",
x"08002FDD",
x"20030000",
x"E8600003",
x"44000806",
x"08002FE1",
x"47A00801",
x"EAC10003",
x"44200006",
x"08002FE5",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"08002FF8",
x"44000806",
x"44210002",
x"47600802",
x"E7E10238",
x"46200001",
x"47600002",
x"E7E00234",
x"08003196",
x"20040003",
x"48640095",
x"C7E1021C",
x"8DC3FFEC",
x"C4600000",
x"44200801",
x"C7E20214",
x"C460FFF8",
x"44400001",
x"44210802",
x"44000002",
x"44200000",
x"44000004",
x"20030034",
x"C4610000",
x"44010003",
x"E4200000",
x"40210008",
x"C0000051",
x"20210008",
x"44000806",
x"C4200000",
x"44010001",
x"441E0002",
x"46C01001",
x"200300F0",
x"C4630000",
x"200300EC",
x"C4640000",
x"E8500003",
x"44400806",
x"08003020",
x"44400807",
x"EBA10027",
x"E8300003",
x"44200006",
x"08003046",
x"443D0800",
x"EBA10013",
x"E8300003",
x"44200006",
x"08003037",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08003032",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003037",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003046",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08003041",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003046",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003069",
x"443D0801",
x"EBA10013",
x"E8300003",
x"44200006",
x"0800305A",
x"443D0800",
x"EBA10009",
x"E8300003",
x"44200006",
x"08003055",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"0800305A",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003069",
x"443D0801",
x"EBA10009",
x"E8300003",
x"44200006",
x"08003064",
x"443D0800",
x"40210008",
x"C0000DE4",
x"20210008",
x"08003069",
x"443D0801",
x"40210008",
x"C0000DE4",
x"20210008",
x"E8600006",
x"EA020003",
x"20030000",
x"0800306E",
x"20030001",
x"08003073",
x"EA020003",
x"20030001",
x"08003073",
x"20030000",
x"E8600003",
x"44000806",
x"08003077",
x"47A00801",
x"EAC10003",
x"44200006",
x"0800307B",
x"44610001",
x"44150802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44800802",
x"44000002",
x"46200000",
x"44200003",
x"48600003",
x"44000807",
x"0800308E",
x"44000806",
x"44210002",
x"441B0802",
x"E7E10234",
x"46200001",
x"441B0002",
x"E7E00230",
x"08003196",
x"20040004",
x"48640100",
x"C7E1021C",
x"8DC5FFEC",
x"C4A00000",
x"44200801",
x"8DC6FFF0",
x"C4C00000",
x"44000004",
x"44200802",
x"C7E20214",
x"C4A0FFF8",
x"44401001",
x"C4C0FFF8",
x"44000004",
x"44401002",
x"44211802",
x"44420002",
x"44602800",
x"E8300003",
x"44200006",
x"080030AC",
x"44200007",
x"2003008C",
x"C4660000",
x"E806005D",
x"44410803",
x"E8300003",
x"44200006",
x"080030B4",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"080030B9",
x"2003FFFF",
x"080030BB",
x"20030001",
x"48600003",
x"44002006",
x"080030BF",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44610803",
x"47201002",
x"47410800",
x"44411003",
x"2004004C",
x"C4810000",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800803",
x"68030006",
x"68600003",
x"44200006",
x"08003104",
x"47E10001",
x"08003106",
x"46C10001",
x"20030044",
x"C4610000",
x"44010002",
x"441E0003",
x"0800310D",
x"20030088",
x"C4600000",
x"E4200004",
x"4021000C",
x"C0000051",
x"2021000C",
x"44000806",
x"C4200004",
x"44013801",
x"C7E10218",
x"C4A0FFFC",
x"44200801",
x"C4C0FFFC",
x"44000004",
x"44200802",
x"E8B00003",
x"44A00006",
x"0800311E",
x"44A00007",
x"E806005D",
x"44250803",
x"E8300003",
x"44200006",
x"08003124",
x"44200007",
x"EA200006",
x"E8140003",
x"20030000",
x"08003129",
x"2003FFFF",
x"0800312B",
x"20030001",
x"48600003",
x"44002006",
x"0800312F",
x"46202003",
x"44840002",
x"20040084",
x"C4810000",
x"44201002",
x"20040080",
x"C4810000",
x"44411003",
x"2004007C",
x"C4810000",
x"44201802",
x"20040078",
x"C4810000",
x"44220800",
x"44611003",
x"20040074",
x"C4810000",
x"44201802",
x"20040070",
x"C4810000",
x"44220800",
x"44611003",
x"2004006C",
x"C4810000",
x"44201802",
x"20040068",
x"C4810000",
x"44220800",
x"44611003",
x"20040064",
x"C4810000",
x"44201802",
x"47820800",
x"44611003",
x"20040060",
x"C4810000",
x"44201802",
x"2004005C",
x"C4810000",
x"44220800",
x"44611003",
x"20040058",
x"C4810000",
x"44201802",
x"20040054",
x"C4810000",
x"44220800",
x"44611003",
x"20040050",
x"C4810000",
x"44201802",
x"47220800",
x"44611003",
x"47200802",
x"47421000",
x"44220803",
x"2004004C",
x"C4820000",
x"44401002",
x"47010800",
x"44410803",
x"46E10800",
x"44010003",
x"46200000",
x"44800003",
x"68030006",
x"68600003",
x"44000806",
x"08003174",
x"47E00801",
x"08003176",
x"46C00801",
x"20030044",
x"C4600000",
x"44200002",
x"441E0003",
x"0800317D",
x"20030088",
x"C4600000",
x"E4200008",
x"40210010",
x"C0000051",
x"20210010",
x"44000806",
x"C4200008",
x"44010001",
x"2003003C",
x"C4620000",
x"46A70801",
x"44210802",
x"44410801",
x"46A00001",
x"44000002",
x"44200801",
x"E8300003",
x"44200006",
x"08003190",
x"46000006",
x"47600802",
x"20030038",
x"C4600000",
x"44200003",
x"E7E00230",
x"08003196",
x"200C0000",
x"8FED0204",
x"40210010",
x"C0002162",
x"20210010",
x"48600025",
x"C7E1022C",
x"C7E00134",
x"44201002",
x"C7E10228",
x"C7E00130",
x"44200002",
x"44401000",
x"C7E10224",
x"C7E0012C",
x"44200002",
x"44400800",
x"44200807",
x"EA010003",
x"46000006",
x"080031AC",
x"44200006",
x"45400802",
x"8DC3FFE4",
x"C4600000",
x"44200002",
x"C7E20244",
x"C7E10238",
x"44010802",
x"44410800",
x"E7E10244",
x"C7E20240",
x"C7E10234",
x"44010802",
x"44410800",
x"E7E10240",
x"C7E2023C",
x"C7E10230",
x"44010002",
x"44400000",
x"E7E0023C",
x"E0000000",
x"E0000000",
x"6B200090",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"080031E3",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"43390002",
x"6B20006C",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"08003206",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"43390002",
x"6B200048",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"08003229",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"43390002",
x"6B200024",
x"A3230002",
x"4EE31800",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E810000A",
x"A3230002",
x"4EE32000",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"0800324C",
x"23230001",
x"A0630002",
x"4EE32000",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210004",
x"C0002EC2",
x"20210004",
x"43390002",
x"080031C1",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"20030004",
x"687A03E8",
x"A3430002",
x"4DA31800",
x"686003E4",
x"A3430002",
x"4D831800",
x"AC390000",
x"AC290004",
x"AC2A0008",
x"AC2B000C",
x"AC2C0010",
x"AC2D0014",
x"AC2E0018",
x"AC2F001C",
x"48600002",
x"08003630",
x"A3430002",
x"4D431800",
x"C4600000",
x"E7E00244",
x"C460FFFC",
x"E7E00240",
x"C460FFF8",
x"E7E0023C",
x"8D3E0000",
x"A3430002",
x"4F23B000",
x"A3430002",
x"4DC3C000",
x"AC2B0020",
x"AC360024",
x"AC380028",
x"4BC00002",
x"0800332C",
x"8FF702CC",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"080032CA",
x"20050002",
x"68A60002",
x"080032CA",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"080032C4",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"080032C9",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C0001DDC",
x"20210030",
x"080032D0",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080032ED",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"0800330A",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"08003327",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00031C1",
x"20210030",
x"4BDC0002",
x"080033E7",
x"8FF702C8",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08003384",
x"20050002",
x"68A60002",
x"08003384",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"0800337E",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"08003383",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C0001DDC",
x"20210030",
x"0800338A",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080033A8",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080033C5",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080033E2",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00031C1",
x"20210030",
x"20030002",
x"4BC30002",
x"080034A3",
x"8FF702C4",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"08003440",
x"20050002",
x"68A60002",
x"08003440",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"0800343A",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"0800343F",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C0001DDC",
x"20210030",
x"08003446",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"08003464",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"08003481",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"0800349E",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00031C1",
x"20210030",
x"20030003",
x"4BC30002",
x"0800355F",
x"8FF702C0",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"080034FC",
x"20050002",
x"68A60002",
x"080034FC",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"080034F6",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"080034FB",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C0001DDC",
x"20210030",
x"08003502",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"08003520",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"0800353D",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"0800355A",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"20030070",
x"20790000",
x"40210030",
x"C00031C1",
x"20210030",
x"20030004",
x"4BC30002",
x"0800361B",
x"8FF702BC",
x"8C380028",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40630001",
x"68600052",
x"A0640002",
x"03E42020",
x"8C840110",
x"8C87FFD8",
x"8C86FFFC",
x"C7010000",
x"8C85FFEC",
x"C4A00000",
x"44200001",
x"E4E00000",
x"C701FFFC",
x"C4A0FFFC",
x"44200001",
x"E4E0FFFC",
x"C701FFF8",
x"C4A0FFF8",
x"44200001",
x"E4E0FFF8",
x"20050002",
x"48C5000F",
x"8C84FFF0",
x"C4E10000",
x"C4E3FFFC",
x"C4E2FFF8",
x"C4800000",
x"44010802",
x"C480FFFC",
x"44030002",
x"44200800",
x"C480FFF8",
x"44020002",
x"44200000",
x"E4E0FFF4",
x"080035B8",
x"20050002",
x"68A60002",
x"080035B8",
x"C4E20000",
x"C4E1FFFC",
x"C4E0FFF8",
x"44422002",
x"8C85FFF0",
x"C4A30000",
x"44832802",
x"44212002",
x"C4A3FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C4A3FFF8",
x"44831802",
x"44A32000",
x"8C85FFF4",
x"48A00003",
x"44801806",
x"080035B2",
x"44202802",
x"8C84FFDC",
x"C4830000",
x"44A31802",
x"44832000",
x"44021802",
x"C480FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C480FFF8",
x"44201802",
x"44831800",
x"20040003",
x"48C40003",
x"44710001",
x"080035B7",
x"44600006",
x"E4E0FFF4",
x"40640001",
x"23030000",
x"40210030",
x"C0001DDC",
x"20210030",
x"080035BE",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"8C360024",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080035DC",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"080035F9",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"08003616",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210030",
x"C0002EC2",
x"20210030",
x"201E0070",
x"23D90000",
x"40210030",
x"C00031C1",
x"20210030",
x"A3430002",
x"8C2B0020",
x"4D631800",
x"C7E20250",
x"C4610000",
x"C7E00244",
x"44200002",
x"44400000",
x"E7E00250",
x"C7E2024C",
x"C461FFFC",
x"C7E00240",
x"44200002",
x"44400000",
x"E7E0024C",
x"C7E20248",
x"C461FFF8",
x"C7E0023C",
x"44200002",
x"44400000",
x"E7E00248",
x"235A0001",
x"8C2F001C",
x"8C2E0018",
x"8C2D0014",
x"8C2C0010",
x"8C2B000C",
x"8C2A0008",
x"8C290004",
x"8C390000",
x"08003252",
x"E0000000",
x"E0000000",
x"A0830002",
x"4CA33000",
x"20030004",
x"687A00A0",
x"8CC7FFF8",
x"A3430002",
x"4CE31800",
x"6860009B",
x"A0870002",
x"4D273800",
x"8CECFFF8",
x"A34B0002",
x"4D8B5800",
x"4963001D",
x"A08B0002",
x"4D0B5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"49630015",
x"408B0001",
x"A16B0002",
x"4CAB5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"4963000C",
x"208B0001",
x"A16B0002",
x"4CAB5800",
x"8D6CFFF8",
x"A34B0002",
x"4D8B5800",
x"49630003",
x"200B0001",
x"08003661",
x"200B0000",
x"08003663",
x"200B0000",
x"08003665",
x"200B0000",
x"08003667",
x"200B0000",
x"4960000C",
x"A0830002",
x"4CA31800",
x"8C79FFE4",
x"8C69FFE8",
x"8C6AFFEC",
x"8C6BFFF0",
x"8C6CFFF4",
x"8C6DFFF8",
x"8C6EFFFC",
x"8C6F0000",
x"08003252",
x"8CCBFFF4",
x"A3430002",
x"4D631800",
x"48600002",
x"080036DC",
x"8CE7FFEC",
x"40830001",
x"A0630002",
x"4CA31800",
x"8C6BFFEC",
x"8CC6FFEC",
x"20830001",
x"A0630002",
x"4CA31800",
x"8C6CFFEC",
x"A0830002",
x"4D031800",
x"8C6DFFEC",
x"A3430002",
x"4CE31800",
x"C4600000",
x"E7E00244",
x"C460FFFC",
x"E7E00240",
x"C460FFF8",
x"E7E0023C",
x"A3430002",
x"4D631800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4CC31800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4D831800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A3430002",
x"4DA31800",
x"C7E10244",
x"C4600000",
x"44200000",
x"E7E00244",
x"C7E10240",
x"C460FFFC",
x"44200000",
x"E7E00240",
x"C7E1023C",
x"C460FFF8",
x"44200000",
x"E7E0023C",
x"A0830002",
x"4CA31800",
x"8C66FFF0",
x"A3430002",
x"4CC31800",
x"C7E20250",
x"C4610000",
x"C7E00244",
x"44200002",
x"44400000",
x"E7E00250",
x"C7E2024C",
x"C461FFFC",
x"C7E00240",
x"44200002",
x"44400000",
x"E7E0024C",
x"C7E20248",
x"C461FFF8",
x"C7E0023C",
x"44200002",
x"44400000",
x"E7E00248",
x"235A0001",
x"0800363C",
x"E0000000",
x"E0000000",
x"20030004",
x"687A00E2",
x"A3430002",
x"4D631800",
x"686000DE",
x"A3430002",
x"4D431800",
x"AC390000",
x"AC2D0004",
x"AC2A0008",
x"AC2B000C",
x"AC2C0010",
x"AC2E0014",
x"48600002",
x"080037BA",
x"8F230000",
x"E7F00244",
x"E7F00240",
x"E7F0023C",
x"A0630002",
x"03E31820",
x"8C7702CC",
x"A3430002",
x"4FC3B000",
x"A3430002",
x"4D83C000",
x"C7000000",
x"E7E0027C",
x"C700FFFC",
x"E7E00278",
x"C700FFF8",
x"E7E00274",
x"8FE3001C",
x"40670001",
x"68E00052",
x"A0E30002",
x"03E31820",
x"8C630110",
x"8C66FFD8",
x"8C65FFFC",
x"C7010000",
x"8C64FFEC",
x"C4800000",
x"44200001",
x"E4C00000",
x"C701FFFC",
x"C480FFFC",
x"44200001",
x"E4C0FFFC",
x"C701FFF8",
x"C480FFF8",
x"44200001",
x"E4C0FFF8",
x"20040002",
x"48A4000F",
x"8C63FFF0",
x"C4C10000",
x"C4C3FFFC",
x"C4C2FFF8",
x"C4600000",
x"44010802",
x"C460FFFC",
x"44030002",
x"44200800",
x"C460FFF8",
x"44020002",
x"44200000",
x"E4C0FFF4",
x"0800374E",
x"20040002",
x"68850002",
x"0800374E",
x"C4C20000",
x"C4C1FFFC",
x"C4C0FFF8",
x"44422002",
x"8C64FFF0",
x"C4830000",
x"44832802",
x"44212002",
x"C483FFFC",
x"44831802",
x"44A32800",
x"44002002",
x"C483FFF8",
x"44831802",
x"44A32000",
x"8C64FFF4",
x"48800003",
x"44801806",
x"08003748",
x"44202802",
x"8C63FFDC",
x"C4630000",
x"44A31802",
x"44832000",
x"44021802",
x"C460FFFC",
x"44600002",
x"44802000",
x"44410802",
x"C460FFF8",
x"44201802",
x"44831800",
x"20030003",
x"48A30003",
x"44710001",
x"0800374D",
x"44600006",
x"E4C0FFF4",
x"40E40001",
x"23030000",
x"4021001C",
x"C0001DDC",
x"2021001C",
x"08003754",
x"8EE3FE28",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"AC290018",
x"E8100009",
x"8EE4FE28",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"08003772",
x"8EE4FE24",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"8EE3FE30",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE30",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"0800378F",
x"8EE4FE2C",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"8EE3FE38",
x"8C630000",
x"C4610000",
x"C6C00000",
x"44201002",
x"C461FFFC",
x"C6C0FFFC",
x"44200002",
x"44401000",
x"C461FFF8",
x"C6C0FFF8",
x"44200002",
x"44400000",
x"E8100009",
x"8EE4FE38",
x"44125003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"080037AC",
x"8EE4FE34",
x"44135003",
x"8C83FFFC",
x"8C950000",
x"40210020",
x"C0002EC2",
x"20210020",
x"20030070",
x"20790000",
x"40210020",
x"C00031C1",
x"20210020",
x"8C290018",
x"A3430002",
x"4D231800",
x"C7E00244",
x"E4600000",
x"C7E00240",
x"E460FFFC",
x"C7E0023C",
x"E460FFF8",
x"235A0001",
x"8C2E0014",
x"8C2C0010",
x"8C2B000C",
x"8C2A0008",
x"8C2D0004",
x"8C390000",
x"080036E0",
x"E0000000",
x"E0000000",
x"68C00076",
x"C7E30264",
x"8FE30260",
x"00C31822",
x"40210004",
x"C0000081",
x"20210004",
x"44600002",
x"C7E10288",
x"44010802",
x"442D0800",
x"E7E102AC",
x"C7E10284",
x"44010802",
x"442C0800",
x"E7E102A8",
x"C7E10280",
x"44010002",
x"440B0000",
x"E7E002A4",
x"C7E202AC",
x"44420802",
x"C7E002A8",
x"44000002",
x"44200800",
x"C7E002A4",
x"44000002",
x"44200000",
x"44000004",
x"C8100003",
x"46200803",
x"080037E6",
x"200300C8",
x"C4610000",
x"44410002",
x"E7E002AC",
x"C7E002A8",
x"44010002",
x"E7E002A8",
x"C7E002A4",
x"44010002",
x"E7E002A4",
x"E7F00250",
x"E7F0024C",
x"E7F00248",
x"C7E00128",
x"E7E00270",
x"C7E00124",
x"E7E0026C",
x"C7E00120",
x"E7E00268",
x"20190000",
x"A0C30002",
x"4CE31800",
x"8C70FFE4",
x"8C75FFE8",
x"8C77FFEC",
x"8C71FFF0",
x"8C72FFF4",
x"8C73FFF8",
x"8C74FFFC",
x"8C780000",
x"43F602AC",
x"E42B0000",
x"E42C0004",
x"E42D0008",
x"AC28000C",
x"AC270010",
x"AC260014",
x"46007006",
x"46206806",
x"4021001C",
x"C0002AAB",
x"2021001C",
x"8C260014",
x"A0C30002",
x"8C270010",
x"4CE31800",
x"8C630000",
x"C7E00250",
x"E4600000",
x"C7E0024C",
x"E460FFFC",
x"C7E00248",
x"E460FFF8",
x"A0C30002",
x"4CE31800",
x"8C63FFE8",
x"8C28000C",
x"AC680000",
x"A0C30002",
x"4CE31800",
x"201A0000",
x"8C7EFFE4",
x"8C79FFE8",
x"8C69FFEC",
x"8C6DFFF0",
x"8C6AFFF4",
x"8C6BFFF8",
x"8C6CFFFC",
x"8C6E0000",
x"4021001C",
x"C00036E0",
x"2021001C",
x"8C260014",
x"40C60001",
x"8C28000C",
x"21030001",
x"20080005",
x"68680003",
x"40680005",
x"08003835",
x"20680000",
x"C42D0008",
x"C42C0004",
x"C42B0000",
x"8C270010",
x"080037C4",
x"E0000000",
x"8FE30258",
x"69C30002",
x"E0000000",
x"A1C30002",
x"4E031800",
x"8C630000",
x"C4600000",
x"E7E00250",
x"C460FFFC",
x"E7E0024C",
x"C460FFF8",
x"E7E00248",
x"8FE40254",
x"21E30001",
x"68640003",
x"20030000",
x"08003858",
x"680F0003",
x"20030000",
x"08003858",
x"8FE40258",
x"21C30001",
x"68640003",
x"20030000",
x"08003858",
x"680E0003",
x"20030000",
x"08003858",
x"20030001",
x"AC320000",
x"AC300004",
x"AC310008",
x"AC2F000C",
x"AC2E0010",
x"48600012",
x"A1C30002",
x"4E032000",
x"201A0000",
x"8C99FFE4",
x"8C89FFE8",
x"8C8AFFEC",
x"8C8BFFF0",
x"8C8CFFF4",
x"8C8DFFF8",
x"8C83FFFC",
x"8C840000",
x"206E0000",
x"208F0000",
x"40210018",
x"C0003252",
x"20210018",
x"08003878",
x"201A0000",
x"22480000",
x"22050000",
x"22290000",
x"21EA0000",
x"21C40000",
x"40210018",
x"C000363C",
x"20210018",
x"C7E00250",
x"40210018",
x"C00000A0",
x"20210018",
x"200400FF",
x"68830006",
x"68600003",
x"20640000",
x"08003882",
x"20040000",
x"08003884",
x"200400FF",
x"40210018",
x"C0001037",
x"20030020",
x"04600001",
x"C7E0024C",
x"C00000A0",
x"20210018",
x"200400FF",
x"68830006",
x"68600003",
x"20640000",
x"08003891",
x"20040000",
x"08003893",
x"200400FF",
x"40210018",
x"C0001037",
x"20030020",
x"04600001",
x"C7E00248",
x"C00000A0",
x"20210018",
x"200400FF",
x"68830006",
x"68600003",
x"20640000",
x"080038A0",
x"20040000",
x"080038A2",
x"200400FF",
x"40210018",
x"C0001037",
x"20210018",
x"2003000A",
x"04600001",
x"8C2E0010",
x"21CE0001",
x"8C2F000C",
x"8C310008",
x"8C300004",
x"8C320000",
x"0800383B",
x"8FE30254",
x"69E30002",
x"E0000000",
x"40630001",
x"AC280000",
x"AC300004",
x"AC310008",
x"AC27000C",
x"AC2F0010",
x"69E30002",
x"080038D1",
x"21E40001",
x"C7E30264",
x"8FE3025C",
x"00831822",
x"40210018",
x"C0000081",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"22070000",
x"C00037C4",
x"20210018",
x"200E0000",
x"8C2F0010",
x"8C27000C",
x"8C310008",
x"8C300004",
x"22120000",
x"22300000",
x"20F10000",
x"40210018",
x"C000383B",
x"20210018",
x"8C2F0010",
x"21EF0001",
x"8C280000",
x"21030002",
x"20080005",
x"68680003",
x"40680005",
x"080038E5",
x"20680000",
x"8FE30254",
x"69E30002",
x"E0000000",
x"40630001",
x"AC280014",
x"AC2F0018",
x"69E30002",
x"08003907",
x"21E40001",
x"C7E30264",
x"8FE3025C",
x"00831822",
x"40210020",
x"C0000081",
x"20210020",
x"44600002",
x"C7E10294",
x"44011002",
x"C7E102A0",
x"44416800",
x"C7E10290",
x"44011002",
x"C7E1029C",
x"44416000",
x"C7E1028C",
x"44010802",
x"C7E00298",
x"44205800",
x"8FE30258",
x"40660001",
x"8C27000C",
x"40210020",
x"C00037C4",
x"20210020",
x"200E0000",
x"8C2F0018",
x"8C310008",
x"8C300004",
x"8C27000C",
x"20F20000",
x"40210020",
x"C000383B",
x"20210020",
x"8C2F0018",
x"21EF0001",
x"8C280014",
x"21040002",
x"20030005",
x"68830003",
x"40830005",
x"08003919",
x"20830000",
x"8C300004",
x"8C27000C",
x"8C310008",
x"20680000",
x"221B0000",
x"22300000",
x"20F10000",
x"23670000",
x"080038AE",
x"6920007D",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"206D0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20680000",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"AD03FFF0",
x"20030005",
x"20040000",
x"C000003F",
x"206C0000",
x"20030005",
x"20040000",
x"C000003F",
x"206B0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20670000",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"ACE3FFF0",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20660000",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"ACC3FFF0",
x"20030001",
x"20040000",
x"C000003F",
x"206E0000",
x"20030003",
x"46000006",
x"C0000048",
x"20640000",
x"20030005",
x"C000003F",
x"20650000",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFFC",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFF8",
x"20030003",
x"46000006",
x"C0000048",
x"ACA3FFF4",
x"20030003",
x"46000006",
x"C0000048",
x"20210004",
x"ACA3FFF0",
x"20430000",
x"20420020",
x"AC65FFE4",
x"AC6EFFE8",
x"AC66FFEC",
x"AC67FFF0",
x"AC6BFFF4",
x"AC6CFFF8",
x"AC68FFFC",
x"AC6D0000",
x"A1240002",
x"6D441800",
x"41290001",
x"08003922",
x"21430000",
x"E0000000",
x"E4200000",
x"E4220004",
x"20060005",
x"68860039",
x"44A51002",
x"44210002",
x"44400000",
x"44110000",
x"44000004",
x"44A01003",
x"44200803",
x"46200003",
x"A0A40002",
x"03E42020",
x"8C8502CC",
x"A0640002",
x"4CA42000",
x"8C840000",
x"E4820000",
x"E481FFFC",
x"E480FFF8",
x"20640028",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44202007",
x"E4820000",
x"E480FFFC",
x"E484FFF8",
x"20640050",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44401807",
x"E4800000",
x"E483FFFC",
x"E484FFF8",
x"20640001",
x"A0840002",
x"4CA42000",
x"8C840000",
x"44000007",
x"E4830000",
x"E484FFFC",
x"E480FFF8",
x"20640029",
x"A0840002",
x"4CA42000",
x"8C840000",
x"E4830000",
x"E480FFFC",
x"E481FFF8",
x"20630051",
x"A0630002",
x"4CA31800",
x"8C630000",
x"E4600000",
x"E462FFFC",
x"E461FFF8",
x"E0000000",
x"44210002",
x"200600A4",
x"C4C60000",
x"44060000",
x"44002804",
x"46250003",
x"EA200006",
x"E8140003",
x"20060000",
x"080039E8",
x"2006FFFF",
x"080039EA",
x"20060001",
x"48C00003",
x"44002006",
x"080039EE",
x"46202003",
x"44840002",
x"20070084",
x"C4EE0000",
x"45C00802",
x"20070080",
x"C4EF0000",
x"442F1803",
x"2007007C",
x"C4E10000",
x"E4210008",
x"C4210008",
x"44201002",
x"20070078",
x"C4E10000",
x"E421000C",
x"C421000C",
x"44230800",
x"44410803",
x"20070074",
x"C4EB0000",
x"45601002",
x"20070070",
x"C4ED0000",
x"45A10800",
x"44411003",
x"2007006C",
x"C4EC0000",
x"45801802",
x"20070068",
x"C4E10000",
x"E4210010",
x"C4210010",
x"44220800",
x"44610803",
x"20070064",
x"C4E90000",
x"45201002",
x"47810800",
x"44411003",
x"20070060",
x"C4EA0000",
x"45401802",
x"2007005C",
x"C4E10000",
x"E4210014",
x"C4210014",
x"44220800",
x"44611003",
x"2007004C",
x"C4E10000",
x"E4210018",
x"20070058",
x"C4E80000",
x"45001802",
x"20070054",
x"C4E10000",
x"E421001C",
x"C421001C",
x"44220800",
x"44610803",
x"20070050",
x"C4E70000",
x"44E01002",
x"47210800",
x"44410803",
x"47201002",
x"47410800",
x"44411003",
x"C4210018",
x"44201802",
x"47020800",
x"44610803",
x"46E10800",
x"44010003",
x"46200000",
x"44800803",
x"68060006",
x"68C00003",
x"44200006",
x"08003A3F",
x"47E10001",
x"08003A41",
x"46C10001",
x"C4210004",
x"44010802",
x"44210002",
x"44191003",
x"47421001",
x"44021003",
x"47021001",
x"44021003",
x"46E21001",
x"44020003",
x"46200001",
x"44200003",
x"44052802",
x"20840001",
x"44A50002",
x"44060000",
x"44003004",
x"46260003",
x"EA200006",
x"E8140003",
x"20060000",
x"08003A58",
x"2006FFFF",
x"08003A5A",
x"20060001",
x"48C00003",
x"44000806",
x"08003A5E",
x"46200803",
x"44210002",
x"45C01002",
x"444F1803",
x"C4220008",
x"44402002",
x"C422000C",
x"44431000",
x"44821003",
x"45601802",
x"45A21000",
x"44621803",
x"45802002",
x"C4220010",
x"44431000",
x"44821003",
x"45201802",
x"47821000",
x"44621003",
x"45401802",
x"C4240014",
x"44821000",
x"44621003",
x"45002002",
x"C423001C",
x"44621000",
x"44821003",
x"44E01802",
x"47221000",
x"44621003",
x"47201802",
x"47421000",
x"44621003",
x"C4230018",
x"44601802",
x"47021000",
x"44621003",
x"46E21000",
x"44020003",
x"46200000",
x"44200803",
x"68060006",
x"68C00003",
x"44200006",
x"08003A8B",
x"47E10001",
x"08003A8D",
x"46C10001",
x"C4210000",
x"44010002",
x"44001002",
x"44590803",
x"47410801",
x"44410803",
x"47010801",
x"44410803",
x"46E10801",
x"44410803",
x"46210801",
x"44010003",
x"44060802",
x"C4220004",
x"C4200000",
x"080039A1",
x"694000AA",
x"E4200000",
x"21430000",
x"40210008",
x"C0000081",
x"20210008",
x"44000806",
x"200300AC",
x"C4650000",
x"44250802",
x"200300A8",
x"C4640000",
x"44241001",
x"20040000",
x"C4200000",
x"E4240004",
x"E4250008",
x"E421000C",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210014",
x"C00039A1",
x"20210014",
x"200300A4",
x"C4630000",
x"C421000C",
x"44231000",
x"20040000",
x"210B0002",
x"C4200000",
x"E4230010",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210018",
x"C00039A1",
x"20210018",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003ACC",
x"20690000",
x"6940007A",
x"21430000",
x"40210018",
x"C0000081",
x"20210018",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E4210014",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"4021001C",
x"C00039A1",
x"2021001C",
x"C4230010",
x"C4210014",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"4021001C",
x"C00039A1",
x"2021001C",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003AF3",
x"20690000",
x"69400052",
x"21430000",
x"4021001C",
x"C0000081",
x"2021001C",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E4210018",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210020",
x"C00039A1",
x"20210020",
x"C4230010",
x"C4210018",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210020",
x"C00039A1",
x"20210020",
x"414A0001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003B1A",
x"20690000",
x"6940002A",
x"21430000",
x"40210020",
x"C0000081",
x"20210020",
x"44000806",
x"C4250008",
x"44250802",
x"C4240004",
x"44241001",
x"20040000",
x"C4200000",
x"E421001C",
x"21030000",
x"21250000",
x"46000806",
x"46002806",
x"40210024",
x"C00039A1",
x"20210024",
x"C4230010",
x"C421001C",
x"44231000",
x"20040000",
x"C4200000",
x"21630000",
x"21250000",
x"46000806",
x"46002806",
x"40210024",
x"C00039A1",
x"20210024",
x"414A0001",
x"21240001",
x"20030005",
x"68830003",
x"40830005",
x"08003B41",
x"20830000",
x"C4200000",
x"20690000",
x"08003A9D",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"69A00132",
x"21A30000",
x"40210004",
x"C0000081",
x"20210004",
x"200300AC",
x"C4640000",
x"44040002",
x"200300A8",
x"C4630000",
x"44030001",
x"20030004",
x"E4200000",
x"40210008",
x"C0000081",
x"20210008",
x"44000806",
x"44240802",
x"44235001",
x"20040000",
x"C4200000",
x"E42A0004",
x"E4230008",
x"E424000C",
x"E4210010",
x"21030000",
x"21850000",
x"45401006",
x"46000806",
x"46002806",
x"40210018",
x"C00039A1",
x"20210018",
x"200300A4",
x"C4650000",
x"C4210010",
x"44254800",
x"20040000",
x"210A0002",
x"C4200000",
x"E4290014",
x"E4250018",
x"21430000",
x"21850000",
x"45201006",
x"46000806",
x"46002806",
x"40210020",
x"C00039A1",
x"20210020",
x"20060003",
x"21830001",
x"20090005",
x"68690003",
x"40690005",
x"08003B81",
x"20690000",
x"20C30000",
x"40210020",
x"C0000081",
x"20210020",
x"44000806",
x"C424000C",
x"44240802",
x"C4230008",
x"44234001",
x"20040000",
x"C4200000",
x"E428001C",
x"E4210020",
x"21030000",
x"21250000",
x"45001006",
x"46000806",
x"46002806",
x"40210028",
x"C00039A1",
x"20210028",
x"C4250018",
x"C4210020",
x"44253800",
x"20040000",
x"C4200000",
x"E4270024",
x"21430000",
x"21250000",
x"44E01006",
x"46000806",
x"46002806",
x"4021002C",
x"C00039A1",
x"2021002C",
x"20060002",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003BAB",
x"20690000",
x"20C30000",
x"4021002C",
x"C0000081",
x"2021002C",
x"44000806",
x"C424000C",
x"44240802",
x"C4230008",
x"44233001",
x"20040000",
x"C4200000",
x"E4260028",
x"E421002C",
x"21030000",
x"21250000",
x"44C01006",
x"46000806",
x"46002806",
x"40210034",
x"C00039A1",
x"20210034",
x"C4250018",
x"C421002C",
x"44251000",
x"20040000",
x"C4200000",
x"E4220030",
x"21430000",
x"21250000",
x"46000806",
x"46002806",
x"40210038",
x"C00039A1",
x"20210038",
x"20060001",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003BD4",
x"20690000",
x"20C30000",
x"40210038",
x"C0000081",
x"20210038",
x"44000806",
x"C424000C",
x"44245802",
x"C4230008",
x"45630801",
x"20040000",
x"C4200000",
x"E42B0034",
x"21030000",
x"21250000",
x"44201006",
x"46002806",
x"46000806",
x"4021003C",
x"C00039A1",
x"2021003C",
x"C4250018",
x"C42B0034",
x"45650800",
x"20040000",
x"C4200000",
x"21430000",
x"21250000",
x"44201006",
x"46002806",
x"46000806",
x"4021003C",
x"C00039A1",
x"2021003C",
x"200A0000",
x"21230001",
x"20090005",
x"68690003",
x"40690005",
x"08003BFC",
x"20690000",
x"C4200000",
x"AC280038",
x"40210040",
x"C0003A9D",
x"20210040",
x"41AE0001",
x"21830002",
x"200C0005",
x"686C0003",
x"406C0005",
x"08003C08",
x"206C0000",
x"8C280038",
x"210D0004",
x"69C0006F",
x"21C30000",
x"40210040",
x"C0000081",
x"20210040",
x"C424000C",
x"44040002",
x"C4230008",
x"44030001",
x"20040000",
x"C42A0004",
x"E420003C",
x"21A30000",
x"21850000",
x"45401006",
x"46000806",
x"46002806",
x"40210044",
x"C00039A1",
x"20210044",
x"20040000",
x"21A80002",
x"C4290014",
x"C420003C",
x"21030000",
x"21850000",
x"45201006",
x"46000806",
x"46002806",
x"40210044",
x"C00039A1",
x"20210044",
x"21830001",
x"20050005",
x"68650003",
x"40650005",
x"08003C30",
x"20650000",
x"20040000",
x"C428001C",
x"C420003C",
x"AC250040",
x"21A30000",
x"45001006",
x"46000806",
x"46002806",
x"40210048",
x"C00039A1",
x"20210048",
x"20040000",
x"C4270024",
x"C420003C",
x"8C250040",
x"21030000",
x"44E01006",
x"46000806",
x"46002806",
x"40210048",
x"C00039A1",
x"20210048",
x"8C250040",
x"20A30001",
x"20050005",
x"68650003",
x"40650005",
x"08003C4D",
x"20650000",
x"20040000",
x"C4260028",
x"C420003C",
x"AC250044",
x"21A30000",
x"44C01006",
x"46000806",
x"46002806",
x"4021004C",
x"C00039A1",
x"2021004C",
x"20040000",
x"C4220030",
x"C420003C",
x"8C250044",
x"21030000",
x"46000806",
x"46002806",
x"4021004C",
x"C00039A1",
x"2021004C",
x"200A0001",
x"8C250044",
x"20A30001",
x"20090005",
x"68690003",
x"40690005",
x"08003C6A",
x"20690000",
x"C420003C",
x"21A80000",
x"4021004C",
x"C0003A9D",
x"2021004C",
x"41C40001",
x"21830002",
x"200C0005",
x"686C0003",
x"406C0005",
x"08003C76",
x"206C0000",
x"21A80004",
x"208D0000",
x"08003B48",
x"E0000000",
x"E0000000",
x"68E00058",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20640000",
x"8FE3001C",
x"AC240000",
x"40210008",
x"C000003F",
x"20210008",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240000",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E00042",
x"20030003",
x"46000006",
x"40210008",
x"C0000048",
x"20210008",
x"20640000",
x"8FE3001C",
x"AC240004",
x"4021000C",
x"C000003F",
x"2021000C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240004",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E0002C",
x"20030003",
x"46000006",
x"4021000C",
x"C0000048",
x"2021000C",
x"20640000",
x"8FE3001C",
x"AC240008",
x"40210010",
x"C000003F",
x"20210010",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240008",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"68E00016",
x"20030003",
x"46000006",
x"40210010",
x"C0000048",
x"20210010",
x"20640000",
x"8FE3001C",
x"AC24000C",
x"40210014",
x"C000003F",
x"20210014",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24000C",
x"AC640000",
x"A0E40002",
x"6CC41800",
x"40E70001",
x"08003C7B",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"690000C2",
x"20060078",
x"20030003",
x"46000006",
x"40210004",
x"C0000048",
x"20210004",
x"20640000",
x"8FE3001C",
x"AC240000",
x"40210008",
x"C000003F",
x"20210008",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240000",
x"AC640000",
x"20640000",
x"20C30000",
x"40210008",
x"C000003F",
x"A1040002",
x"03E42020",
x"AC8302CC",
x"A1030002",
x"03E31820",
x"8C6602CC",
x"20030003",
x"46000006",
x"C0000048",
x"20210008",
x"20640000",
x"8FE3001C",
x"AC240004",
x"4021000C",
x"C000003F",
x"2021000C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240004",
x"AC640000",
x"ACC3FE28",
x"20030003",
x"46000006",
x"4021000C",
x"C0000048",
x"2021000C",
x"20640000",
x"8FE3001C",
x"AC240008",
x"40210010",
x"C000003F",
x"20210010",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240008",
x"AC640000",
x"ACC3FE2C",
x"20030003",
x"46000006",
x"40210010",
x"C0000048",
x"20210010",
x"20640000",
x"8FE3001C",
x"AC24000C",
x"40210014",
x"C000003F",
x"20210014",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24000C",
x"AC640000",
x"ACC3FE30",
x"20030003",
x"46000006",
x"40210014",
x"C0000048",
x"20210014",
x"20640000",
x"8FE3001C",
x"AC240010",
x"40210018",
x"C000003F",
x"20210018",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240010",
x"AC640000",
x"ACC3FE34",
x"20070072",
x"40210018",
x"C0003C7B",
x"20210018",
x"41080001",
x"69000058",
x"20060078",
x"20030003",
x"46000006",
x"40210018",
x"C0000048",
x"20210018",
x"20640000",
x"8FE3001C",
x"AC240014",
x"4021001C",
x"C000003F",
x"2021001C",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240014",
x"AC640000",
x"20640000",
x"20C30000",
x"4021001C",
x"C000003F",
x"A1040002",
x"03E42020",
x"AC8302CC",
x"A1030002",
x"03E31820",
x"8C6602CC",
x"20030003",
x"46000006",
x"C0000048",
x"2021001C",
x"20640000",
x"8FE3001C",
x"AC240018",
x"40210020",
x"C000003F",
x"20210020",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240018",
x"AC640000",
x"ACC3FE28",
x"20030003",
x"46000006",
x"40210020",
x"C0000048",
x"20210020",
x"20640000",
x"8FE3001C",
x"AC24001C",
x"40210024",
x"C000003F",
x"20210024",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C24001C",
x"AC640000",
x"ACC3FE2C",
x"20030003",
x"46000006",
x"40210024",
x"C0000048",
x"20210024",
x"20640000",
x"8FE3001C",
x"AC240020",
x"40210028",
x"C000003F",
x"20210028",
x"20650000",
x"20430000",
x"20420008",
x"AC65FFFC",
x"8C240020",
x"AC640000",
x"ACC3FE30",
x"20070073",
x"40210028",
x"C0003C7B",
x"20210028",
x"41080001",
x"08003CD4",
x"E0000000",
x"E0000000",
x"69800060",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"69800054",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"69800048",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"6980003C",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"69800030",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"69800024",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"69800018",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"6980000C",
x"A1830002",
x"4D631800",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"20210004",
x"418C0001",
x"08003D97",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"E0000000",
x"69A0006E",
x"A1A30002",
x"03E31820",
x"8C6B02CC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE40",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"200C006F",
x"C0003D97",
x"20210004",
x"41AD0001",
x"69A00034",
x"A1A30002",
x"03E31820",
x"8C6B02CC",
x"8D63FE24",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"40210004",
x"C0001D15",
x"8D63FE28",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE2C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE30",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE34",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE38",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"8D63FE3C",
x"8FE4001C",
x"40850001",
x"8C66FFFC",
x"8C670000",
x"C0001D15",
x"200C0070",
x"C0003D97",
x"20210004",
x"41AD0001",
x"08003DF8",
x"E0000000",
x"E0000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000"

	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



