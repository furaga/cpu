library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
--use ieee.std_logic_signed.all;

entity prom is
	port (
		clka : in std_logic;
		addra : in std_logic_vector(9 downto 0);
		douta : out std_logic_vector(31 downto 0));



end prom;

architecture RTL of prom is
	subtype word_t is std_logic_vector(31 downto 0);
	type mem_t is array (0 to 1023) of word_t;
	signal addr_in	: integer range 0 to 1023;

	constant mem : mem_t := (
x"0000004C",
x"00000000",
x"3F800000",
x"BF800000",
x"00800000",
x"4B000000",
x"4B000000",
x"41400000",
x"41300000",
x"41200000",
x"41100000",
x"41000000",
x"40E00000",
x"40C00000",
x"40A00000",
x"40800000",
x"40400000",
x"3F800000",
x"00000000",
x"40000000",
x"08000098",
x"A0630002",
x"00622820",
x"20430000",
x"68A20005",
x"28A20004",
x"AC440000",
x"20420004",
x"08000018",
x"E0000000",
x"A0630002",
x"00622020",
x"20430000",
x"68820005",
x"28820004",
x"E4400000",
x"20420004",
x"08000021",
x"E0000000",
x"44000806",
x"20030000",
x"C4640000",
x"E8800015",
x"C8800014",
x"44000007",
x"20030010",
x"C4620000",
x"E8020004",
x"C8020003",
x"44000007",
x"E0000000",
x"44020000",
x"44020001",
x"44200807",
x"E820001B",
x"C820001A",
x"44020000",
x"20030004",
x"C4630000",
x"44030000",
x"44020001",
x"44000007",
x"E0000000",
x"20030010",
x"C4620000",
x"E8020003",
x"C8020002",
x"E0000000",
x"44000806",
x"44020000",
x"E4200000",
x"8C240000",
x"44020001",
x"E4200000",
x"8C240000",
x"E8010005",
x"C8010004",
x"20030004",
x"C4630000",
x"44030001",
x"E0000000",
x"44000007",
x"E0000000",
x"44000007",
x"C0000027",
x"44000007",
x"E0000000",
x"68030006",
x"28030005",
x"00031822",
x"C000005D",
x"44000007",
x"E0000000",
x"20050010",
x"C4A10000",
x"20050014",
x"8CA40000",
x"2005000C",
x"8CA50000",
x"68A30007",
x"28A30006",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"E0000000",
x"20040000",
x"C4820000",
x"00651822",
x"44411000",
x"68A3FFFE",
x"28A3FFFD",
x"00641820",
x"AC230000",
x"C4200000",
x"44010001",
x"44020000",
x"E0000000",
x"20030000",
x"C4610000",
x"E8200006",
x"C8200005",
x"44000007",
x"C000007E",
x"00031822",
x"E0000000",
x"C0000027",
x"20040010",
x"C4820000",
x"20040014",
x"8C840000",
x"E8400007",
x"C8400006",
x"44020000",
x"E4200000",
x"8C230000",
x"00641822",
x"E0000000",
x"2005000C",
x"8CA50000",
x"20030000",
x"44020001",
x"00651820",
x"E840FFFE",
x"C840FFFD",
x"44020000",
x"E4200000",
x"8C250000",
x"00A42822",
x"00A31820",
x"E0000000",
x"08000076",
x"203F0000",
x"40210030",
x"201C0001",
x"201DFFFF",
x"201B0044",
x"C7700000",
x"201B0020",
x"C7710000",
x"201B0024",
x"C7720000",
x"201B0028",
x"C7730000",
x"201B002C",
x"C7740000",
x"201B0030",
x"C7750000",
x"201B0034",
x"C7760000",
x"201B0038",
x"C7770000",
x"201B003C",
x"C7780000",
x"201B0040",
x"C7790000",
x"201B0048",
x"C77A0000",
x"201B0018",
x"C77B0000",
x"201B001C",
x"C77C0000",
x"47400006",
x"20030001",
x"20040000",
x"AFE2002C",
x"43E20004",
x"E4200000",
x"40210008",
x"C0000015",
x"8FE2002C",
x"20030001",
x"20040000",
x"AFE2002C",
x"43E20008",
x"C0000015",
x"8FE2002C",
x"20030001",
x"20040000",
x"AFE2002C",
x"43E2000C",
x"C0000015",
x"8FE2002C",
x"20030001",
x"20040000",
x"AFE2002C",
x"43E20010",
x"C0000015",
x"8FE2002C",
x"20030001",
x"20040001",
x"AFE2002C",
x"43E20014",
x"C0000015",
x"8FE2002C",
x"20030001",
x"20040000",
x"AFE2002C",
x"43E20018",
x"C0000015",
x"8FE2002C",
x"20030000",
x"46000006",
x"AFE2002C",
x"43E2001C",
x"C000001E",
x"8FE2002C",
x"20030002",
x"20040003",
x"C00002C2",
x"20210008",
x"AFE30020",
x"20040003",
x"20050002",
x"AC230004",
x"20830000",
x"20A40000",
x"4021000C",
x"C00002C2",
x"2021000C",
x"AFE30024",
x"20040002",
x"20050002",
x"AC230008",
x"20830000",
x"20A40000",
x"40210010",
x"C00002C2",
x"20210010",
x"20680000",
x"AFE80028",
x"8C260004",
x"8CC30000",
x"47200006",
x"E4600000",
x"8CC30000",
x"C4200000",
x"E460FFFC",
x"8CC30000",
x"47000006",
x"E460FFF8",
x"8CC3FFFC",
x"46E00006",
x"E4600000",
x"8CC3FFFC",
x"46C00006",
x"E460FFFC",
x"8CC3FFFC",
x"46A00006",
x"E460FFF8",
x"8C270008",
x"8CE30000",
x"46800006",
x"E4600000",
x"8CE30000",
x"46600006",
x"E460FFFC",
x"8CE3FFFC",
x"46400006",
x"E4600000",
x"8CE3FFFC",
x"46200006",
x"E460FFFC",
x"8CE3FFF8",
x"47800006",
x"E4600000",
x"8CE3FFF8",
x"47600006",
x"E460FFFC",
x"20030002",
x"20040003",
x"20050002",
x"AC28000C",
x"40210014",
x"C00002A2",
x"20210014",
x"8C23000C",
x"8C640000",
x"C4800000",
x"40210014",
x"C0000097",
x"C0000164",
x"20210014",
x"AC230014",
x"2003000A",
x"04600001",
x"8C230014",
x"8C23000C",
x"8C640000",
x"C480FFFC",
x"40210014",
x"C0000097",
x"C0000164",
x"20210014",
x"AC230014",
x"2003000A",
x"04600001",
x"8C230014",
x"8C23000C",
x"8C64FFFC",
x"C4800000",
x"40210014",
x"C0000097",
x"C0000164",
x"20210014",
x"AC230014",
x"2003000A",
x"04600001",
x"8C230014",
x"8C23000C",
x"8C63FFFC",
x"C460FFFC",
x"40210014",
x"C0000097",
x"C0000164",
x"20210014",
x"AC230014",
x"2003000A",
x"04600001",
x"8C230014",
x"0000003F",
x"00A63820",
x"A8E70001",
x"00E44018",
x"00C54822",
x"6B890003",
x"20A30000",
x"E0000000",
x"69030006",
x"49030003",
x"20E30000",
x"E0000000",
x"20E60000",
x"08000155",
x"20E50000",
x"08000155",
x"686000E2",
x"3C8005F5",
x"1C80E100",
x"20050000",
x"20060003",
x"AC230000",
x"40210008",
x"C0000155",
x"20210008",
x"3C8005F5",
x"1C80E100",
x"00642018",
x"8C250000",
x"00A42022",
x"AC240004",
x"68030003",
x"20030000",
x"0800017A",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"3C800098",
x"1C809680",
x"20050000",
x"2006000A",
x"8C270004",
x"AC230008",
x"20E30000",
x"40210010",
x"C0000155",
x"20210010",
x"3C800098",
x"1C809680",
x"00642018",
x"8C250004",
x"00A42022",
x"AC24000C",
x"6803000A",
x"8C250008",
x"48A00003",
x"20030000",
x"08000193",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"08000198",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"3C80000F",
x"1C804240",
x"20050000",
x"2006000A",
x"8C27000C",
x"AC230010",
x"20E30000",
x"40210018",
x"C0000155",
x"20210018",
x"3C80000F",
x"1C804240",
x"00642018",
x"8C25000C",
x"00A42022",
x"AC240014",
x"6803000A",
x"8C250010",
x"48A00003",
x"20030000",
x"080001B1",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"080001B6",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"3C800001",
x"1C8086A0",
x"20050000",
x"2006000A",
x"8C270014",
x"AC230018",
x"20E30000",
x"40210020",
x"C0000155",
x"20210020",
x"3C800001",
x"1C8086A0",
x"00642018",
x"8C250014",
x"00A42022",
x"AC24001C",
x"6803000A",
x"8C250018",
x"48A00003",
x"20030000",
x"080001CF",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"080001D4",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"20042710",
x"20050000",
x"2006000A",
x"8C27001C",
x"AC230020",
x"20E30000",
x"40210028",
x"C0000155",
x"20210028",
x"20042710",
x"00642018",
x"8C25001C",
x"00A42022",
x"AC240024",
x"6803000A",
x"8C250020",
x"48A00003",
x"20030000",
x"080001EB",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"080001F0",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"200403E8",
x"20050000",
x"2006000A",
x"8C270024",
x"AC230028",
x"20E30000",
x"40210030",
x"C0000155",
x"20210030",
x"606403E8",
x"8C250024",
x"00A42022",
x"AC24002C",
x"6803000A",
x"8C250028",
x"48A00003",
x"20030000",
x"08000206",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"0800020B",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"20040064",
x"20050000",
x"2006000A",
x"8C27002C",
x"AC230030",
x"20E30000",
x"40210038",
x"C0000155",
x"20210038",
x"60640064",
x"8C25002C",
x"00A42022",
x"AC240034",
x"6803000A",
x"8C250030",
x"48A00003",
x"20030000",
x"08000221",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"08000226",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"2004000A",
x"20050000",
x"2006000A",
x"8C270034",
x"AC230038",
x"20E30000",
x"40210040",
x"C0000155",
x"20210040",
x"6064000A",
x"8C250034",
x"00A42022",
x"AC24003C",
x"6803000A",
x"8C250038",
x"48A00003",
x"20030000",
x"0800023C",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"08000241",
x"20050030",
x"00A31820",
x"04600001",
x"20030001",
x"20030030",
x"8C24003C",
x"00641820",
x"04600001",
x"E0000000",
x"2004002D",
x"AC230000",
x"04800001",
x"8C230000",
x"00031822",
x"08000164",
x"8FC4FFEC",
x"8FC5FFF0",
x"8FC6FFF4",
x"8FC7FFF8",
x"8FC8FFFC",
x"68600014",
x"A0A90002",
x"4CC93000",
x"A0890002",
x"00C90031",
x"A0A50002",
x"4D052800",
x"A0680002",
x"00A80831",
x"A0650002",
x"4CE52800",
x"A0870002",
x"00A71031",
x"44220802",
x"44010000",
x"A0840002",
x"00C40039",
x"40630001",
x"8FDB0000",
x"03600008",
x"E0000000",
x"8FC4FFEC",
x"8FC5FFF0",
x"8FC6FFF4",
x"8FC7FFF8",
x"8FC8FFFC",
x"68600018",
x"20490000",
x"20420018",
x"200A024C",
x"AD2A0000",
x"AD23FFEC",
x"AD25FFF0",
x"AD26FFF4",
x"AD27FFF8",
x"AD28FFFC",
x"40840001",
x"AC3E0000",
x"AC230004",
x"20830000",
x"213E0000",
x"8FDB0000",
x"4021000C",
x"03600030",
x"2021000C",
x"8C230004",
x"40630001",
x"8C3E0000",
x"8FDB0000",
x"03600008",
x"E0000000",
x"8FC4FFEC",
x"8FC5FFF0",
x"8FC6FFF4",
x"8FC7FFF8",
x"8FC8FFFC",
x"68600018",
x"20490000",
x"20420018",
x"200A0266",
x"AD2A0000",
x"AD25FFEC",
x"AD23FFF0",
x"AD26FFF4",
x"AD27FFF8",
x"AD28FFFC",
x"40840001",
x"AC3E0000",
x"AC230004",
x"20830000",
x"213E0000",
x"8FDB0000",
x"4021000C",
x"03600030",
x"2021000C",
x"8C230004",
x"40630001",
x"8C3E0000",
x"8FDB0000",
x"03600008",
x"E0000000",
x"205E0000",
x"20420018",
x"20090284",
x"AFC90000",
x"AFC5FFEC",
x"AFC4FFF0",
x"AFC8FFF4",
x"AFC7FFF8",
x"AFC6FFFC",
x"40630001",
x"8FDB0000",
x"03600008",
x"8FC4FFF8",
x"8FC5FFFC",
x"68600011",
x"46000006",
x"AC3E0000",
x"AC250004",
x"AC230008",
x"20830000",
x"40210010",
x"C000001E",
x"20210010",
x"8C240008",
x"A0850002",
x"8C260004",
x"6CC51800",
x"40830001",
x"8C3E0000",
x"8FDB0000",
x"03600008",
x"E0000000",
x"43E5001C",
x"AC230000",
x"AC240004",
x"20A40000",
x"4021000C",
x"C0000015",
x"2021000C",
x"205E0000",
x"2042000C",
x"200402AE",
x"AFC40000",
x"8C240004",
x"AFC4FFF8",
x"AFC3FFFC",
x"8C240000",
x"40840001",
x"AC230008",
x"20830000",
x"8FDB0000",
x"40210010",
x"03600030",
x"20210010",
x"8C230008",
x"E0000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000"

	 );


begin
	prom_sim: process(clka)
	begin
		if rising_edge(clka) then
			addr_in <= conv_integer(addra);
			douta <= mem(addr_in);
		end if;
	end process;

end RTL;



